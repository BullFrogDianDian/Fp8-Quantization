module ControlUnit(
  input  [31:0] io_addr, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  input  [31:0] io_data, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output        io_encoderLinearConfig_en, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output        io_encoderLinearConfig_weight, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_encoderLinearConfig_i, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_encoderLinearConfig_j, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_encoderLinearConfig_value, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output        io_decoderLinearConfig_en, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output        io_decoderLinearConfig_weight, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_decoderLinearConfig_i, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_decoderLinearConfig_j, // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
  output [7:0]  io_decoderLinearConfig_value // @[src/main/scala/Multiple/ControlUnit.scala 18:20]
);
  wire [11:0] cs = io_addr[27:16]; // @[src/main/scala/Multiple/ControlUnit.scala 25:25]
  wire  _T = cs == 12'h1; // @[src/main/scala/Multiple/ControlUnit.scala 32:18]
  wire  _T_2 = cs == 12'h3; // @[src/main/scala/Multiple/ControlUnit.scala 46:17]
  assign io_encoderLinearConfig_en = cs == 12'h2 | _T; // @[src/main/scala/Multiple/ControlUnit.scala 36:31 37:43]
  assign io_encoderLinearConfig_weight = cs == 12'h2 ? 1'h0 : 1'h1; // @[src/main/scala/Multiple/ControlUnit.scala 36:31 38:47]
  assign io_encoderLinearConfig_i = io_addr[15:8]; // @[src/main/scala/Multiple/ControlUnit.scala 29:44]
  assign io_encoderLinearConfig_j = io_addr[7:0]; // @[src/main/scala/Multiple/ControlUnit.scala 30:44]
  assign io_encoderLinearConfig_value = io_data[7:0]; // @[src/main/scala/Multiple/ControlUnit.scala 31:48]
  assign io_decoderLinearConfig_en = cs == 12'h4 | _T_2; // @[src/main/scala/Multiple/ControlUnit.scala 50:30 51:43]
  assign io_decoderLinearConfig_weight = cs == 12'h4 ? 1'h0 : 1'h1; // @[src/main/scala/Multiple/ControlUnit.scala 50:30 52:47]
  assign io_decoderLinearConfig_i = io_addr[15:8]; // @[src/main/scala/Multiple/ControlUnit.scala 43:44]
  assign io_decoderLinearConfig_j = io_addr[7:0]; // @[src/main/scala/Multiple/ControlUnit.scala 44:44]
  assign io_decoderLinearConfig_value = io_data[7:0]; // @[src/main/scala/Multiple/ControlUnit.scala 45:48]
endmodule
module LinearCompute(
  input           clock,
  input           io_pipe_validIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output          io_pipe_validOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_en, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_weight, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_i, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_j, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_value, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_63, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_31, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_scale, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_zeroPoint // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [2047:0] _RAND_9;
  reg [2047:0] _RAND_10;
  reg [2047:0] _RAND_11;
  reg [2047:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] linear_weight_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [31:0] ansAll_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [31:0] ansAll_63_0_extendedIn1 = {24'h0,io_featuresIn_63}; // @[src/main/scala/Multiple/LinearCompute.scala 29:30]
  wire [31:0] ansAll_63_31_extendedIn2 = {24'h0,linear_weight_63_31}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_63_31_product = ansAll_63_0_extendedIn1 * ansAll_63_31_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  reg [7:0] ans_31; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [31:0] tempSum_31; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  wire [31:0] _GEN_10336 = {{16'd0}, io_zeroPoint}; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] biasExtended_31 = {24'h0,linear_bias_31}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_31 = tempSum_31 + biasExtended_31; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_31_sign = sum32_31[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_31_absX_T = ~sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_31_absX_T_2 = _ans_31_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_31_absX = ans_31_sign ? _ans_31_absX_T_2 : sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_31_shiftedX_T_1 = _GEN_10336 - ans_31_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_31_shiftedX_T_3 = ans_31_absX - _GEN_10336; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_31_shiftedX = ans_31_sign ? _ans_31_shiftedX_T_1 : _ans_31_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_31_scaledX_T_1 = ans_31_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_31_scaledX = _ans_31_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_31_clippedX_T_2 = ans_31_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_31_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_31_clippedX = ans_31_scaledX > 49'h1c0 ? 49'h1c0 : _ans_31_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_31_absClipped_T_1 = ~ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_31_absClipped_T_3 = _ans_31_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_31_absClipped = ans_31_clippedX[31] ? _ans_31_absClipped_T_3 : ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_31_isZero = ans_31_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10679 = {{16'd0}, ans_31_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_4 = _GEN_10679 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_6 = {ans_31_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_8 = _ans_31_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_9 = _ans_31_leadingZeros_T_4 | _ans_31_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10680 = {{8'd0}, _ans_31_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_14 = _GEN_10680 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_16 = {_ans_31_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_18 = _ans_31_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_19 = _ans_31_leadingZeros_T_14 | _ans_31_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10681 = {{4'd0}, _ans_31_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_24 = _GEN_10681 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_26 = {_ans_31_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_28 = _ans_31_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_29 = _ans_31_leadingZeros_T_24 | _ans_31_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10682 = {{2'd0}, _ans_31_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_34 = _GEN_10682 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_36 = {_ans_31_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_38 = _ans_31_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_39 = _ans_31_leadingZeros_T_34 | _ans_31_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10683 = {{1'd0}, _ans_31_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_44 = _GEN_10683 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_46 = {_ans_31_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_48 = _ans_31_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_49 = _ans_31_leadingZeros_T_44 | _ans_31_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10684 = {{8'd0}, ans_31_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_55 = _GEN_10684 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_57 = {ans_31_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_59 = _ans_31_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_60 = _ans_31_leadingZeros_T_55 | _ans_31_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10685 = {{4'd0}, _ans_31_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_65 = _GEN_10685 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_67 = {_ans_31_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_69 = _ans_31_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_70 = _ans_31_leadingZeros_T_65 | _ans_31_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10686 = {{2'd0}, _ans_31_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_75 = _GEN_10686 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_77 = {_ans_31_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_79 = _ans_31_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_80 = _ans_31_leadingZeros_T_75 | _ans_31_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10687 = {{1'd0}, _ans_31_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_85 = _GEN_10687 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_87 = {_ans_31_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_89 = _ans_31_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_90 = _ans_31_leadingZeros_T_85 | _ans_31_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_31_leadingZeros_T_93 = {_ans_31_leadingZeros_T_49,_ans_31_leadingZeros_T_90,ans_31_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_31_leadingZeros_T_143 = _ans_31_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_144 = _ans_31_leadingZeros_T_93[46] ? 6'h2e : _ans_31_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_145 = _ans_31_leadingZeros_T_93[45] ? 6'h2d : _ans_31_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_146 = _ans_31_leadingZeros_T_93[44] ? 6'h2c : _ans_31_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_147 = _ans_31_leadingZeros_T_93[43] ? 6'h2b : _ans_31_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_148 = _ans_31_leadingZeros_T_93[42] ? 6'h2a : _ans_31_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_149 = _ans_31_leadingZeros_T_93[41] ? 6'h29 : _ans_31_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_150 = _ans_31_leadingZeros_T_93[40] ? 6'h28 : _ans_31_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_151 = _ans_31_leadingZeros_T_93[39] ? 6'h27 : _ans_31_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_152 = _ans_31_leadingZeros_T_93[38] ? 6'h26 : _ans_31_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_153 = _ans_31_leadingZeros_T_93[37] ? 6'h25 : _ans_31_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_154 = _ans_31_leadingZeros_T_93[36] ? 6'h24 : _ans_31_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_155 = _ans_31_leadingZeros_T_93[35] ? 6'h23 : _ans_31_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_156 = _ans_31_leadingZeros_T_93[34] ? 6'h22 : _ans_31_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_157 = _ans_31_leadingZeros_T_93[33] ? 6'h21 : _ans_31_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_158 = _ans_31_leadingZeros_T_93[32] ? 6'h20 : _ans_31_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_159 = _ans_31_leadingZeros_T_93[31] ? 6'h1f : _ans_31_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_160 = _ans_31_leadingZeros_T_93[30] ? 6'h1e : _ans_31_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_161 = _ans_31_leadingZeros_T_93[29] ? 6'h1d : _ans_31_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_162 = _ans_31_leadingZeros_T_93[28] ? 6'h1c : _ans_31_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_163 = _ans_31_leadingZeros_T_93[27] ? 6'h1b : _ans_31_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_164 = _ans_31_leadingZeros_T_93[26] ? 6'h1a : _ans_31_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_165 = _ans_31_leadingZeros_T_93[25] ? 6'h19 : _ans_31_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_166 = _ans_31_leadingZeros_T_93[24] ? 6'h18 : _ans_31_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_167 = _ans_31_leadingZeros_T_93[23] ? 6'h17 : _ans_31_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_168 = _ans_31_leadingZeros_T_93[22] ? 6'h16 : _ans_31_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_169 = _ans_31_leadingZeros_T_93[21] ? 6'h15 : _ans_31_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_170 = _ans_31_leadingZeros_T_93[20] ? 6'h14 : _ans_31_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_171 = _ans_31_leadingZeros_T_93[19] ? 6'h13 : _ans_31_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_172 = _ans_31_leadingZeros_T_93[18] ? 6'h12 : _ans_31_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_173 = _ans_31_leadingZeros_T_93[17] ? 6'h11 : _ans_31_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_174 = _ans_31_leadingZeros_T_93[16] ? 6'h10 : _ans_31_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_175 = _ans_31_leadingZeros_T_93[15] ? 6'hf : _ans_31_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_176 = _ans_31_leadingZeros_T_93[14] ? 6'he : _ans_31_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_177 = _ans_31_leadingZeros_T_93[13] ? 6'hd : _ans_31_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_178 = _ans_31_leadingZeros_T_93[12] ? 6'hc : _ans_31_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_179 = _ans_31_leadingZeros_T_93[11] ? 6'hb : _ans_31_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_180 = _ans_31_leadingZeros_T_93[10] ? 6'ha : _ans_31_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_181 = _ans_31_leadingZeros_T_93[9] ? 6'h9 : _ans_31_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_182 = _ans_31_leadingZeros_T_93[8] ? 6'h8 : _ans_31_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_183 = _ans_31_leadingZeros_T_93[7] ? 6'h7 : _ans_31_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_184 = _ans_31_leadingZeros_T_93[6] ? 6'h6 : _ans_31_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_185 = _ans_31_leadingZeros_T_93[5] ? 6'h5 : _ans_31_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_186 = _ans_31_leadingZeros_T_93[4] ? 6'h4 : _ans_31_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_187 = _ans_31_leadingZeros_T_93[3] ? 6'h3 : _ans_31_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_188 = _ans_31_leadingZeros_T_93[2] ? 6'h2 : _ans_31_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_189 = _ans_31_leadingZeros_T_93[1] ? 6'h1 : _ans_31_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_31_leadingZeros = _ans_31_leadingZeros_T_93[0] ? 6'h0 : _ans_31_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_expRaw_T_1 = 6'h1f - ans_31_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_31_expRaw = ans_31_isZero ? 6'h0 : _ans_31_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_31_shiftAmt_T_2 = ans_31_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_31_shiftAmt = ans_31_expRaw > 6'h3 ? _ans_31_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_31_mantissaRaw_T = ans_31_absClipped >> ans_31_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_31_mantissaRaw = _ans_31_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_31_mantissa = ans_31_expRaw >= 6'h3 ? ans_31_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_31_expAdjusted = ans_31_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_31_exp_T_4 = ans_31_expAdjusted > 7'hf ? 4'hf : ans_31_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_31_exp = ans_31_isZero ? 4'h0 : _ans_31_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_31_fp8 = {ans_31_clippedX[31],ans_31_exp,ans_31_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [7:0] io_featuresOut_31_scaledX = {{2'd0}, ans_31[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_31_sum = io_featuresOut_31_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_31_minVal = io_featuresOut_31_sum < 8'h40 ? io_featuresOut_31_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  reg  regs__0; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__1; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__2; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__3; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg [2047:0] regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  assign io_pipe_validOut = regs__3; // @[src/main/scala/fpga/Pipeline.scala 46:21]
  assign io_pipe_phvOut = regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 37:21]
  assign io_featuresOut_31 = io_featuresOut_31_minVal > 8'h0 ? io_featuresOut_31_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  always @(posedge clock) begin
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3f == io_config_i[5:0] & 5'h1f == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_63_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    ansAll_63_31 <= ansAll_63_31_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    if (ans_31_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_31 <= 8'h0;
    end else begin
      ans_31 <= ans_31_fp8;
    end
    tempSum_31 <= tempSum_31 + ansAll_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    regs__0 <= io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 45:25]
    regs__1 <= regs__0; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__2 <= regs__1; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__3 <= regs__2; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs_1_0 <= io_pipe_phvIn; // @[src/main/scala/fpga/Pipeline.scala 36:25]
    regs_1_1 <= regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_2 <= regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_3 <= regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 34:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  linear_weight_63_31 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  linear_bias_31 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  ansAll_63_31 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ans_31 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  tempSum_31 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs__0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  regs__1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regs__2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  regs__3 = _RAND_8[0:0];
  _RAND_9 = {64{`RANDOM}};
  regs_1_0 = _RAND_9[2047:0];
  _RAND_10 = {64{`RANDOM}};
  regs_1_1 = _RAND_10[2047:0];
  _RAND_11 = {64{`RANDOM}};
  regs_1_2 = _RAND_11[2047:0];
  _RAND_12 = {64{`RANDOM}};
  regs_1_3 = _RAND_12[2047:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LinearCompute_1(
  input           clock,
  input           io_pipe_validIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output          io_pipe_validOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_en, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_weight, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_i, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_j, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_value, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_31, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_0, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_1, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_2, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_3, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_4, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_5, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_6, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_7, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_8, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_9, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_10, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_11, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_12, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_13, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_14, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_15, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_16, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_17, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_18, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_19, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_20, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_21, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_22, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_23, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_24, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_25, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_26, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_27, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_28, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_29, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_30, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_31, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_32, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_33, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_34, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_35, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_36, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_37, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_38, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_39, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_40, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_41, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_42, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_43, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_44, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_45, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_46, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_47, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_48, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_49, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_50, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_51, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_52, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_53, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_54, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_55, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_56, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_57, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_58, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_59, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_60, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_61, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_62, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_63, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_scale, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_zeroPoint // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [2047:0] _RAND_324;
  reg [2047:0] _RAND_325;
  reg [2047:0] _RAND_326;
  reg [2047:0] _RAND_327;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] linear_weight_31_0; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_1; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_2; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_3; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_4; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_5; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_6; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_7; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_8; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_9; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_10; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_11; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_12; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_13; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_14; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_15; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_16; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_17; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_18; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_19; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_20; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_21; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_22; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_23; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_24; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_25; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_26; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_27; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_28; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_29; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_30; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_32; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_33; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_34; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_35; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_36; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_37; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_38; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_39; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_40; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_41; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_42; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_43; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_44; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_45; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_46; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_47; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_48; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_49; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_50; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_51; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_52; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_53; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_54; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_55; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_56; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_57; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_58; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_59; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_60; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_61; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_62; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_31_63; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_0; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_1; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_2; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_3; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_4; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_5; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_6; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_7; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_8; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_9; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_10; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_11; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_12; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_13; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_14; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_15; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_16; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_17; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_18; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_19; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_20; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_21; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_22; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_23; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_24; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_25; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_26; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_27; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_28; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_29; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_30; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_32; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_33; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_34; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_35; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_36; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_37; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_38; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_39; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_40; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_41; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_42; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_43; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_44; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_45; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_46; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_47; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_48; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_49; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_50; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_51; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_52; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_53; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_54; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_55; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_56; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_57; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_58; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_59; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_60; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_61; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_62; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_63; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [31:0] ansAll_31_0; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_1; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_2; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_3; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_4; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_5; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_6; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_7; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_8; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_9; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_10; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_11; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_12; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_13; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_14; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_15; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_16; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_17; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_18; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_19; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_20; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_21; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_22; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_23; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_24; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_25; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_26; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_27; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_28; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_29; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_30; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_31; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_32; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_33; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_34; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_35; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_36; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_37; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_38; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_39; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_40; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_41; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_42; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_43; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_44; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_45; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_46; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_47; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_48; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_49; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_50; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_51; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_52; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_53; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_54; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_55; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_56; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_57; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_58; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_59; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_60; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_61; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_62; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  reg [31:0] ansAll_31_63; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [31:0] ansAll_31_0_extendedIn1 = {24'h0,io_featuresIn_31}; // @[src/main/scala/Multiple/LinearCompute.scala 29:30]
  wire [31:0] ansAll_31_0_extendedIn2 = {24'h0,linear_weight_31_0}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_0_product = ansAll_31_0_extendedIn1 * ansAll_31_0_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_1_extendedIn2 = {24'h0,linear_weight_31_1}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_1_product = ansAll_31_0_extendedIn1 * ansAll_31_1_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_2_extendedIn2 = {24'h0,linear_weight_31_2}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_2_product = ansAll_31_0_extendedIn1 * ansAll_31_2_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_3_extendedIn2 = {24'h0,linear_weight_31_3}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_3_product = ansAll_31_0_extendedIn1 * ansAll_31_3_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_4_extendedIn2 = {24'h0,linear_weight_31_4}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_4_product = ansAll_31_0_extendedIn1 * ansAll_31_4_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_5_extendedIn2 = {24'h0,linear_weight_31_5}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_5_product = ansAll_31_0_extendedIn1 * ansAll_31_5_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_6_extendedIn2 = {24'h0,linear_weight_31_6}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_6_product = ansAll_31_0_extendedIn1 * ansAll_31_6_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_7_extendedIn2 = {24'h0,linear_weight_31_7}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_7_product = ansAll_31_0_extendedIn1 * ansAll_31_7_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_8_extendedIn2 = {24'h0,linear_weight_31_8}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_8_product = ansAll_31_0_extendedIn1 * ansAll_31_8_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_9_extendedIn2 = {24'h0,linear_weight_31_9}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_9_product = ansAll_31_0_extendedIn1 * ansAll_31_9_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_10_extendedIn2 = {24'h0,linear_weight_31_10}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_10_product = ansAll_31_0_extendedIn1 * ansAll_31_10_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_11_extendedIn2 = {24'h0,linear_weight_31_11}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_11_product = ansAll_31_0_extendedIn1 * ansAll_31_11_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_12_extendedIn2 = {24'h0,linear_weight_31_12}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_12_product = ansAll_31_0_extendedIn1 * ansAll_31_12_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_13_extendedIn2 = {24'h0,linear_weight_31_13}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_13_product = ansAll_31_0_extendedIn1 * ansAll_31_13_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_14_extendedIn2 = {24'h0,linear_weight_31_14}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_14_product = ansAll_31_0_extendedIn1 * ansAll_31_14_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_15_extendedIn2 = {24'h0,linear_weight_31_15}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_15_product = ansAll_31_0_extendedIn1 * ansAll_31_15_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_16_extendedIn2 = {24'h0,linear_weight_31_16}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_16_product = ansAll_31_0_extendedIn1 * ansAll_31_16_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_17_extendedIn2 = {24'h0,linear_weight_31_17}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_17_product = ansAll_31_0_extendedIn1 * ansAll_31_17_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_18_extendedIn2 = {24'h0,linear_weight_31_18}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_18_product = ansAll_31_0_extendedIn1 * ansAll_31_18_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_19_extendedIn2 = {24'h0,linear_weight_31_19}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_19_product = ansAll_31_0_extendedIn1 * ansAll_31_19_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_20_extendedIn2 = {24'h0,linear_weight_31_20}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_20_product = ansAll_31_0_extendedIn1 * ansAll_31_20_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_21_extendedIn2 = {24'h0,linear_weight_31_21}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_21_product = ansAll_31_0_extendedIn1 * ansAll_31_21_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_22_extendedIn2 = {24'h0,linear_weight_31_22}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_22_product = ansAll_31_0_extendedIn1 * ansAll_31_22_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_23_extendedIn2 = {24'h0,linear_weight_31_23}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_23_product = ansAll_31_0_extendedIn1 * ansAll_31_23_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_24_extendedIn2 = {24'h0,linear_weight_31_24}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_24_product = ansAll_31_0_extendedIn1 * ansAll_31_24_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_25_extendedIn2 = {24'h0,linear_weight_31_25}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_25_product = ansAll_31_0_extendedIn1 * ansAll_31_25_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_26_extendedIn2 = {24'h0,linear_weight_31_26}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_26_product = ansAll_31_0_extendedIn1 * ansAll_31_26_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_27_extendedIn2 = {24'h0,linear_weight_31_27}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_27_product = ansAll_31_0_extendedIn1 * ansAll_31_27_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_28_extendedIn2 = {24'h0,linear_weight_31_28}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_28_product = ansAll_31_0_extendedIn1 * ansAll_31_28_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_29_extendedIn2 = {24'h0,linear_weight_31_29}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_29_product = ansAll_31_0_extendedIn1 * ansAll_31_29_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_30_extendedIn2 = {24'h0,linear_weight_31_30}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_30_product = ansAll_31_0_extendedIn1 * ansAll_31_30_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_31_extendedIn2 = {24'h0,linear_weight_31_31}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_31_product = ansAll_31_0_extendedIn1 * ansAll_31_31_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_32_extendedIn2 = {24'h0,linear_weight_31_32}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_32_product = ansAll_31_0_extendedIn1 * ansAll_31_32_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_33_extendedIn2 = {24'h0,linear_weight_31_33}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_33_product = ansAll_31_0_extendedIn1 * ansAll_31_33_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_34_extendedIn2 = {24'h0,linear_weight_31_34}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_34_product = ansAll_31_0_extendedIn1 * ansAll_31_34_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_35_extendedIn2 = {24'h0,linear_weight_31_35}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_35_product = ansAll_31_0_extendedIn1 * ansAll_31_35_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_36_extendedIn2 = {24'h0,linear_weight_31_36}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_36_product = ansAll_31_0_extendedIn1 * ansAll_31_36_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_37_extendedIn2 = {24'h0,linear_weight_31_37}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_37_product = ansAll_31_0_extendedIn1 * ansAll_31_37_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_38_extendedIn2 = {24'h0,linear_weight_31_38}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_38_product = ansAll_31_0_extendedIn1 * ansAll_31_38_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_39_extendedIn2 = {24'h0,linear_weight_31_39}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_39_product = ansAll_31_0_extendedIn1 * ansAll_31_39_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_40_extendedIn2 = {24'h0,linear_weight_31_40}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_40_product = ansAll_31_0_extendedIn1 * ansAll_31_40_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_41_extendedIn2 = {24'h0,linear_weight_31_41}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_41_product = ansAll_31_0_extendedIn1 * ansAll_31_41_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_42_extendedIn2 = {24'h0,linear_weight_31_42}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_42_product = ansAll_31_0_extendedIn1 * ansAll_31_42_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_43_extendedIn2 = {24'h0,linear_weight_31_43}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_43_product = ansAll_31_0_extendedIn1 * ansAll_31_43_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_44_extendedIn2 = {24'h0,linear_weight_31_44}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_44_product = ansAll_31_0_extendedIn1 * ansAll_31_44_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_45_extendedIn2 = {24'h0,linear_weight_31_45}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_45_product = ansAll_31_0_extendedIn1 * ansAll_31_45_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_46_extendedIn2 = {24'h0,linear_weight_31_46}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_46_product = ansAll_31_0_extendedIn1 * ansAll_31_46_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_47_extendedIn2 = {24'h0,linear_weight_31_47}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_47_product = ansAll_31_0_extendedIn1 * ansAll_31_47_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_48_extendedIn2 = {24'h0,linear_weight_31_48}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_48_product = ansAll_31_0_extendedIn1 * ansAll_31_48_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_49_extendedIn2 = {24'h0,linear_weight_31_49}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_49_product = ansAll_31_0_extendedIn1 * ansAll_31_49_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_50_extendedIn2 = {24'h0,linear_weight_31_50}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_50_product = ansAll_31_0_extendedIn1 * ansAll_31_50_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_51_extendedIn2 = {24'h0,linear_weight_31_51}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_51_product = ansAll_31_0_extendedIn1 * ansAll_31_51_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_52_extendedIn2 = {24'h0,linear_weight_31_52}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_52_product = ansAll_31_0_extendedIn1 * ansAll_31_52_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_53_extendedIn2 = {24'h0,linear_weight_31_53}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_53_product = ansAll_31_0_extendedIn1 * ansAll_31_53_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_54_extendedIn2 = {24'h0,linear_weight_31_54}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_54_product = ansAll_31_0_extendedIn1 * ansAll_31_54_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_55_extendedIn2 = {24'h0,linear_weight_31_55}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_55_product = ansAll_31_0_extendedIn1 * ansAll_31_55_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_56_extendedIn2 = {24'h0,linear_weight_31_56}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_56_product = ansAll_31_0_extendedIn1 * ansAll_31_56_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_57_extendedIn2 = {24'h0,linear_weight_31_57}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_57_product = ansAll_31_0_extendedIn1 * ansAll_31_57_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_58_extendedIn2 = {24'h0,linear_weight_31_58}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_58_product = ansAll_31_0_extendedIn1 * ansAll_31_58_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_59_extendedIn2 = {24'h0,linear_weight_31_59}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_59_product = ansAll_31_0_extendedIn1 * ansAll_31_59_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_60_extendedIn2 = {24'h0,linear_weight_31_60}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_60_product = ansAll_31_0_extendedIn1 * ansAll_31_60_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_61_extendedIn2 = {24'h0,linear_weight_31_61}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_61_product = ansAll_31_0_extendedIn1 * ansAll_31_61_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_62_extendedIn2 = {24'h0,linear_weight_31_62}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_62_product = ansAll_31_0_extendedIn1 * ansAll_31_62_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  wire [31:0] ansAll_31_63_extendedIn2 = {24'h0,linear_weight_31_63}; // @[src/main/scala/Multiple/LinearCompute.scala 30:30]
  wire [63:0] ansAll_31_63_product = ansAll_31_0_extendedIn1 * ansAll_31_63_extendedIn2; // @[src/main/scala/Multiple/LinearCompute.scala 31:35]
  reg [7:0] ans_0; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_1; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_2; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_3; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_4; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_5; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_6; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_7; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_8; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_9; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_10; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_11; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_12; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_13; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_14; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_15; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_16; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_17; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_18; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_19; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_20; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_21; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_22; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_23; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_24; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_25; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_26; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_27; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_28; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_29; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_30; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_31; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_32; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_33; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_34; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_35; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_36; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_37; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_38; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_39; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_40; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_41; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_42; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_43; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_44; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_45; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_46; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_47; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_48; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_49; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_50; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_51; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_52; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_53; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_54; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_55; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_56; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_57; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_58; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_59; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_60; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_61; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_62; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [7:0] ans_63; // @[src/main/scala/Multiple/LinearCompute.scala 83:18]
  reg [31:0] tempSum_0; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_1; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_2; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_3; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_4; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_5; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_6; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_7; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_8; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_9; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_10; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_11; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_12; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_13; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_14; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_15; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_16; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_17; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_18; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_19; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_20; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_21; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_22; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_23; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_24; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_25; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_26; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_27; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_28; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_29; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_30; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_31; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_32; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_33; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_34; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_35; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_36; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_37; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_38; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_39; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_40; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_41; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_42; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_43; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_44; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_45; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_46; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_47; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_48; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_49; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_50; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_51; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_52; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_53; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_54; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_55; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_56; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_57; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_58; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_59; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_60; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_61; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_62; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  reg [31:0] tempSum_63; // @[src/main/scala/Multiple/LinearCompute.scala 84:22]
  wire [31:0] biasExtended = {24'h0,linear_bias_0}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32 = tempSum_0 + biasExtended; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_0_sign = sum32[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_0_absX_T = ~sum32; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_0_absX_T_2 = _ans_0_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_0_absX = ans_0_sign ? _ans_0_absX_T_2 : sum32; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _GEN_10432 = {{16'd0}, io_zeroPoint}; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_0_shiftedX_T_1 = _GEN_10432 - ans_0_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_0_shiftedX_T_3 = ans_0_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_0_shiftedX = ans_0_sign ? _ans_0_shiftedX_T_1 : _ans_0_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_0_scaledX_T_1 = ans_0_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_0_scaledX = _ans_0_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_0_clippedX_T_2 = ans_0_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_0_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_0_clippedX = ans_0_scaledX > 49'h1c0 ? 49'h1c0 : _ans_0_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_0_absClipped_T_1 = ~ans_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_0_absClipped_T_3 = _ans_0_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_0_absClipped = ans_0_clippedX[31] ? _ans_0_absClipped_T_3 : ans_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_0_isZero = ans_0_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10434 = {{16'd0}, ans_0_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_4 = _GEN_10434 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_6 = {ans_0_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_8 = _ans_0_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_9 = _ans_0_leadingZeros_T_4 | _ans_0_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10435 = {{8'd0}, _ans_0_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_14 = _GEN_10435 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_16 = {_ans_0_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_18 = _ans_0_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_19 = _ans_0_leadingZeros_T_14 | _ans_0_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10436 = {{4'd0}, _ans_0_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_24 = _GEN_10436 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_26 = {_ans_0_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_28 = _ans_0_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_29 = _ans_0_leadingZeros_T_24 | _ans_0_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10437 = {{2'd0}, _ans_0_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_34 = _GEN_10437 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_36 = {_ans_0_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_38 = _ans_0_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_39 = _ans_0_leadingZeros_T_34 | _ans_0_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10438 = {{1'd0}, _ans_0_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_44 = _GEN_10438 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_46 = {_ans_0_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_48 = _ans_0_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_0_leadingZeros_T_49 = _ans_0_leadingZeros_T_44 | _ans_0_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10439 = {{8'd0}, ans_0_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_55 = _GEN_10439 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_57 = {ans_0_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_59 = _ans_0_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_60 = _ans_0_leadingZeros_T_55 | _ans_0_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10440 = {{4'd0}, _ans_0_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_65 = _GEN_10440 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_67 = {_ans_0_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_69 = _ans_0_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_70 = _ans_0_leadingZeros_T_65 | _ans_0_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10441 = {{2'd0}, _ans_0_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_75 = _GEN_10441 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_77 = {_ans_0_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_79 = _ans_0_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_80 = _ans_0_leadingZeros_T_75 | _ans_0_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10442 = {{1'd0}, _ans_0_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_85 = _GEN_10442 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_87 = {_ans_0_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_89 = _ans_0_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_0_leadingZeros_T_90 = _ans_0_leadingZeros_T_85 | _ans_0_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_0_leadingZeros_T_93 = {_ans_0_leadingZeros_T_49,_ans_0_leadingZeros_T_90,ans_0_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_0_leadingZeros_T_143 = _ans_0_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_144 = _ans_0_leadingZeros_T_93[46] ? 6'h2e : _ans_0_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_145 = _ans_0_leadingZeros_T_93[45] ? 6'h2d : _ans_0_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_146 = _ans_0_leadingZeros_T_93[44] ? 6'h2c : _ans_0_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_147 = _ans_0_leadingZeros_T_93[43] ? 6'h2b : _ans_0_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_148 = _ans_0_leadingZeros_T_93[42] ? 6'h2a : _ans_0_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_149 = _ans_0_leadingZeros_T_93[41] ? 6'h29 : _ans_0_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_150 = _ans_0_leadingZeros_T_93[40] ? 6'h28 : _ans_0_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_151 = _ans_0_leadingZeros_T_93[39] ? 6'h27 : _ans_0_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_152 = _ans_0_leadingZeros_T_93[38] ? 6'h26 : _ans_0_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_153 = _ans_0_leadingZeros_T_93[37] ? 6'h25 : _ans_0_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_154 = _ans_0_leadingZeros_T_93[36] ? 6'h24 : _ans_0_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_155 = _ans_0_leadingZeros_T_93[35] ? 6'h23 : _ans_0_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_156 = _ans_0_leadingZeros_T_93[34] ? 6'h22 : _ans_0_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_157 = _ans_0_leadingZeros_T_93[33] ? 6'h21 : _ans_0_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_158 = _ans_0_leadingZeros_T_93[32] ? 6'h20 : _ans_0_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_159 = _ans_0_leadingZeros_T_93[31] ? 6'h1f : _ans_0_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_160 = _ans_0_leadingZeros_T_93[30] ? 6'h1e : _ans_0_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_161 = _ans_0_leadingZeros_T_93[29] ? 6'h1d : _ans_0_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_162 = _ans_0_leadingZeros_T_93[28] ? 6'h1c : _ans_0_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_163 = _ans_0_leadingZeros_T_93[27] ? 6'h1b : _ans_0_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_164 = _ans_0_leadingZeros_T_93[26] ? 6'h1a : _ans_0_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_165 = _ans_0_leadingZeros_T_93[25] ? 6'h19 : _ans_0_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_166 = _ans_0_leadingZeros_T_93[24] ? 6'h18 : _ans_0_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_167 = _ans_0_leadingZeros_T_93[23] ? 6'h17 : _ans_0_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_168 = _ans_0_leadingZeros_T_93[22] ? 6'h16 : _ans_0_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_169 = _ans_0_leadingZeros_T_93[21] ? 6'h15 : _ans_0_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_170 = _ans_0_leadingZeros_T_93[20] ? 6'h14 : _ans_0_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_171 = _ans_0_leadingZeros_T_93[19] ? 6'h13 : _ans_0_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_172 = _ans_0_leadingZeros_T_93[18] ? 6'h12 : _ans_0_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_173 = _ans_0_leadingZeros_T_93[17] ? 6'h11 : _ans_0_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_174 = _ans_0_leadingZeros_T_93[16] ? 6'h10 : _ans_0_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_175 = _ans_0_leadingZeros_T_93[15] ? 6'hf : _ans_0_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_176 = _ans_0_leadingZeros_T_93[14] ? 6'he : _ans_0_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_177 = _ans_0_leadingZeros_T_93[13] ? 6'hd : _ans_0_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_178 = _ans_0_leadingZeros_T_93[12] ? 6'hc : _ans_0_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_179 = _ans_0_leadingZeros_T_93[11] ? 6'hb : _ans_0_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_180 = _ans_0_leadingZeros_T_93[10] ? 6'ha : _ans_0_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_181 = _ans_0_leadingZeros_T_93[9] ? 6'h9 : _ans_0_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_182 = _ans_0_leadingZeros_T_93[8] ? 6'h8 : _ans_0_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_183 = _ans_0_leadingZeros_T_93[7] ? 6'h7 : _ans_0_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_184 = _ans_0_leadingZeros_T_93[6] ? 6'h6 : _ans_0_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_185 = _ans_0_leadingZeros_T_93[5] ? 6'h5 : _ans_0_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_186 = _ans_0_leadingZeros_T_93[4] ? 6'h4 : _ans_0_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_187 = _ans_0_leadingZeros_T_93[3] ? 6'h3 : _ans_0_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_188 = _ans_0_leadingZeros_T_93[2] ? 6'h2 : _ans_0_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_189 = _ans_0_leadingZeros_T_93[1] ? 6'h1 : _ans_0_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_0_leadingZeros = _ans_0_leadingZeros_T_93[0] ? 6'h0 : _ans_0_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_expRaw_T_1 = 6'h1f - ans_0_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_0_expRaw = ans_0_isZero ? 6'h0 : _ans_0_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_0_shiftAmt_T_2 = ans_0_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_0_shiftAmt = ans_0_expRaw > 6'h3 ? _ans_0_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_0_mantissaRaw_T = ans_0_absClipped >> ans_0_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_0_mantissaRaw = _ans_0_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_0_mantissa = ans_0_expRaw >= 6'h3 ? ans_0_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_0_expAdjusted = ans_0_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_0_exp_T_4 = ans_0_expAdjusted > 7'hf ? 4'hf : ans_0_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_0_exp = ans_0_isZero ? 4'h0 : _ans_0_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_0_fp8 = {ans_0_clippedX[31],ans_0_exp,ans_0_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_1 = {24'h0,linear_bias_1}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_1 = tempSum_1 + biasExtended_1; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_1_sign = sum32_1[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_1_absX_T = ~sum32_1; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_1_absX_T_2 = _ans_1_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_1_absX = ans_1_sign ? _ans_1_absX_T_2 : sum32_1; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_1_shiftedX_T_1 = _GEN_10432 - ans_1_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_1_shiftedX_T_3 = ans_1_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_1_shiftedX = ans_1_sign ? _ans_1_shiftedX_T_1 : _ans_1_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_1_scaledX_T_1 = ans_1_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_1_scaledX = _ans_1_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_1_clippedX_T_2 = ans_1_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_1_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_1_clippedX = ans_1_scaledX > 49'h1c0 ? 49'h1c0 : _ans_1_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_1_absClipped_T_1 = ~ans_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_1_absClipped_T_3 = _ans_1_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_1_absClipped = ans_1_clippedX[31] ? _ans_1_absClipped_T_3 : ans_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_1_isZero = ans_1_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10445 = {{16'd0}, ans_1_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_4 = _GEN_10445 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_6 = {ans_1_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_8 = _ans_1_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_9 = _ans_1_leadingZeros_T_4 | _ans_1_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10446 = {{8'd0}, _ans_1_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_14 = _GEN_10446 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_16 = {_ans_1_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_18 = _ans_1_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_19 = _ans_1_leadingZeros_T_14 | _ans_1_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10447 = {{4'd0}, _ans_1_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_24 = _GEN_10447 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_26 = {_ans_1_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_28 = _ans_1_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_29 = _ans_1_leadingZeros_T_24 | _ans_1_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10448 = {{2'd0}, _ans_1_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_34 = _GEN_10448 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_36 = {_ans_1_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_38 = _ans_1_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_39 = _ans_1_leadingZeros_T_34 | _ans_1_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10449 = {{1'd0}, _ans_1_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_44 = _GEN_10449 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_46 = {_ans_1_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_48 = _ans_1_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_1_leadingZeros_T_49 = _ans_1_leadingZeros_T_44 | _ans_1_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10450 = {{8'd0}, ans_1_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_55 = _GEN_10450 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_57 = {ans_1_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_59 = _ans_1_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_60 = _ans_1_leadingZeros_T_55 | _ans_1_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10451 = {{4'd0}, _ans_1_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_65 = _GEN_10451 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_67 = {_ans_1_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_69 = _ans_1_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_70 = _ans_1_leadingZeros_T_65 | _ans_1_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10452 = {{2'd0}, _ans_1_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_75 = _GEN_10452 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_77 = {_ans_1_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_79 = _ans_1_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_80 = _ans_1_leadingZeros_T_75 | _ans_1_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10453 = {{1'd0}, _ans_1_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_85 = _GEN_10453 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_87 = {_ans_1_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_89 = _ans_1_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_1_leadingZeros_T_90 = _ans_1_leadingZeros_T_85 | _ans_1_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_1_leadingZeros_T_93 = {_ans_1_leadingZeros_T_49,_ans_1_leadingZeros_T_90,ans_1_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_1_leadingZeros_T_143 = _ans_1_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_144 = _ans_1_leadingZeros_T_93[46] ? 6'h2e : _ans_1_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_145 = _ans_1_leadingZeros_T_93[45] ? 6'h2d : _ans_1_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_146 = _ans_1_leadingZeros_T_93[44] ? 6'h2c : _ans_1_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_147 = _ans_1_leadingZeros_T_93[43] ? 6'h2b : _ans_1_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_148 = _ans_1_leadingZeros_T_93[42] ? 6'h2a : _ans_1_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_149 = _ans_1_leadingZeros_T_93[41] ? 6'h29 : _ans_1_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_150 = _ans_1_leadingZeros_T_93[40] ? 6'h28 : _ans_1_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_151 = _ans_1_leadingZeros_T_93[39] ? 6'h27 : _ans_1_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_152 = _ans_1_leadingZeros_T_93[38] ? 6'h26 : _ans_1_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_153 = _ans_1_leadingZeros_T_93[37] ? 6'h25 : _ans_1_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_154 = _ans_1_leadingZeros_T_93[36] ? 6'h24 : _ans_1_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_155 = _ans_1_leadingZeros_T_93[35] ? 6'h23 : _ans_1_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_156 = _ans_1_leadingZeros_T_93[34] ? 6'h22 : _ans_1_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_157 = _ans_1_leadingZeros_T_93[33] ? 6'h21 : _ans_1_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_158 = _ans_1_leadingZeros_T_93[32] ? 6'h20 : _ans_1_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_159 = _ans_1_leadingZeros_T_93[31] ? 6'h1f : _ans_1_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_160 = _ans_1_leadingZeros_T_93[30] ? 6'h1e : _ans_1_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_161 = _ans_1_leadingZeros_T_93[29] ? 6'h1d : _ans_1_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_162 = _ans_1_leadingZeros_T_93[28] ? 6'h1c : _ans_1_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_163 = _ans_1_leadingZeros_T_93[27] ? 6'h1b : _ans_1_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_164 = _ans_1_leadingZeros_T_93[26] ? 6'h1a : _ans_1_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_165 = _ans_1_leadingZeros_T_93[25] ? 6'h19 : _ans_1_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_166 = _ans_1_leadingZeros_T_93[24] ? 6'h18 : _ans_1_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_167 = _ans_1_leadingZeros_T_93[23] ? 6'h17 : _ans_1_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_168 = _ans_1_leadingZeros_T_93[22] ? 6'h16 : _ans_1_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_169 = _ans_1_leadingZeros_T_93[21] ? 6'h15 : _ans_1_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_170 = _ans_1_leadingZeros_T_93[20] ? 6'h14 : _ans_1_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_171 = _ans_1_leadingZeros_T_93[19] ? 6'h13 : _ans_1_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_172 = _ans_1_leadingZeros_T_93[18] ? 6'h12 : _ans_1_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_173 = _ans_1_leadingZeros_T_93[17] ? 6'h11 : _ans_1_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_174 = _ans_1_leadingZeros_T_93[16] ? 6'h10 : _ans_1_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_175 = _ans_1_leadingZeros_T_93[15] ? 6'hf : _ans_1_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_176 = _ans_1_leadingZeros_T_93[14] ? 6'he : _ans_1_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_177 = _ans_1_leadingZeros_T_93[13] ? 6'hd : _ans_1_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_178 = _ans_1_leadingZeros_T_93[12] ? 6'hc : _ans_1_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_179 = _ans_1_leadingZeros_T_93[11] ? 6'hb : _ans_1_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_180 = _ans_1_leadingZeros_T_93[10] ? 6'ha : _ans_1_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_181 = _ans_1_leadingZeros_T_93[9] ? 6'h9 : _ans_1_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_182 = _ans_1_leadingZeros_T_93[8] ? 6'h8 : _ans_1_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_183 = _ans_1_leadingZeros_T_93[7] ? 6'h7 : _ans_1_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_184 = _ans_1_leadingZeros_T_93[6] ? 6'h6 : _ans_1_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_185 = _ans_1_leadingZeros_T_93[5] ? 6'h5 : _ans_1_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_186 = _ans_1_leadingZeros_T_93[4] ? 6'h4 : _ans_1_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_187 = _ans_1_leadingZeros_T_93[3] ? 6'h3 : _ans_1_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_188 = _ans_1_leadingZeros_T_93[2] ? 6'h2 : _ans_1_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_189 = _ans_1_leadingZeros_T_93[1] ? 6'h1 : _ans_1_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_1_leadingZeros = _ans_1_leadingZeros_T_93[0] ? 6'h0 : _ans_1_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_expRaw_T_1 = 6'h1f - ans_1_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_1_expRaw = ans_1_isZero ? 6'h0 : _ans_1_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_1_shiftAmt_T_2 = ans_1_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_1_shiftAmt = ans_1_expRaw > 6'h3 ? _ans_1_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_1_mantissaRaw_T = ans_1_absClipped >> ans_1_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_1_mantissaRaw = _ans_1_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_1_mantissa = ans_1_expRaw >= 6'h3 ? ans_1_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_1_expAdjusted = ans_1_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_1_exp_T_4 = ans_1_expAdjusted > 7'hf ? 4'hf : ans_1_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_1_exp = ans_1_isZero ? 4'h0 : _ans_1_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_1_fp8 = {ans_1_clippedX[31],ans_1_exp,ans_1_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_2 = {24'h0,linear_bias_2}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_2 = tempSum_2 + biasExtended_2; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_2_sign = sum32_2[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_2_absX_T = ~sum32_2; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_2_absX_T_2 = _ans_2_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_2_absX = ans_2_sign ? _ans_2_absX_T_2 : sum32_2; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_2_shiftedX_T_1 = _GEN_10432 - ans_2_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_2_shiftedX_T_3 = ans_2_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_2_shiftedX = ans_2_sign ? _ans_2_shiftedX_T_1 : _ans_2_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_2_scaledX_T_1 = ans_2_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_2_scaledX = _ans_2_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_2_clippedX_T_2 = ans_2_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_2_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_2_clippedX = ans_2_scaledX > 49'h1c0 ? 49'h1c0 : _ans_2_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_2_absClipped_T_1 = ~ans_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_2_absClipped_T_3 = _ans_2_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_2_absClipped = ans_2_clippedX[31] ? _ans_2_absClipped_T_3 : ans_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_2_isZero = ans_2_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10456 = {{16'd0}, ans_2_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_4 = _GEN_10456 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_6 = {ans_2_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_8 = _ans_2_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_9 = _ans_2_leadingZeros_T_4 | _ans_2_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10457 = {{8'd0}, _ans_2_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_14 = _GEN_10457 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_16 = {_ans_2_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_18 = _ans_2_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_19 = _ans_2_leadingZeros_T_14 | _ans_2_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10458 = {{4'd0}, _ans_2_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_24 = _GEN_10458 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_26 = {_ans_2_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_28 = _ans_2_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_29 = _ans_2_leadingZeros_T_24 | _ans_2_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10459 = {{2'd0}, _ans_2_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_34 = _GEN_10459 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_36 = {_ans_2_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_38 = _ans_2_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_39 = _ans_2_leadingZeros_T_34 | _ans_2_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10460 = {{1'd0}, _ans_2_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_44 = _GEN_10460 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_46 = {_ans_2_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_48 = _ans_2_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_2_leadingZeros_T_49 = _ans_2_leadingZeros_T_44 | _ans_2_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10461 = {{8'd0}, ans_2_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_55 = _GEN_10461 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_57 = {ans_2_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_59 = _ans_2_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_60 = _ans_2_leadingZeros_T_55 | _ans_2_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10462 = {{4'd0}, _ans_2_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_65 = _GEN_10462 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_67 = {_ans_2_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_69 = _ans_2_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_70 = _ans_2_leadingZeros_T_65 | _ans_2_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10463 = {{2'd0}, _ans_2_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_75 = _GEN_10463 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_77 = {_ans_2_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_79 = _ans_2_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_80 = _ans_2_leadingZeros_T_75 | _ans_2_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10464 = {{1'd0}, _ans_2_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_85 = _GEN_10464 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_87 = {_ans_2_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_89 = _ans_2_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_2_leadingZeros_T_90 = _ans_2_leadingZeros_T_85 | _ans_2_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_2_leadingZeros_T_93 = {_ans_2_leadingZeros_T_49,_ans_2_leadingZeros_T_90,ans_2_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_2_leadingZeros_T_143 = _ans_2_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_144 = _ans_2_leadingZeros_T_93[46] ? 6'h2e : _ans_2_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_145 = _ans_2_leadingZeros_T_93[45] ? 6'h2d : _ans_2_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_146 = _ans_2_leadingZeros_T_93[44] ? 6'h2c : _ans_2_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_147 = _ans_2_leadingZeros_T_93[43] ? 6'h2b : _ans_2_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_148 = _ans_2_leadingZeros_T_93[42] ? 6'h2a : _ans_2_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_149 = _ans_2_leadingZeros_T_93[41] ? 6'h29 : _ans_2_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_150 = _ans_2_leadingZeros_T_93[40] ? 6'h28 : _ans_2_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_151 = _ans_2_leadingZeros_T_93[39] ? 6'h27 : _ans_2_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_152 = _ans_2_leadingZeros_T_93[38] ? 6'h26 : _ans_2_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_153 = _ans_2_leadingZeros_T_93[37] ? 6'h25 : _ans_2_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_154 = _ans_2_leadingZeros_T_93[36] ? 6'h24 : _ans_2_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_155 = _ans_2_leadingZeros_T_93[35] ? 6'h23 : _ans_2_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_156 = _ans_2_leadingZeros_T_93[34] ? 6'h22 : _ans_2_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_157 = _ans_2_leadingZeros_T_93[33] ? 6'h21 : _ans_2_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_158 = _ans_2_leadingZeros_T_93[32] ? 6'h20 : _ans_2_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_159 = _ans_2_leadingZeros_T_93[31] ? 6'h1f : _ans_2_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_160 = _ans_2_leadingZeros_T_93[30] ? 6'h1e : _ans_2_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_161 = _ans_2_leadingZeros_T_93[29] ? 6'h1d : _ans_2_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_162 = _ans_2_leadingZeros_T_93[28] ? 6'h1c : _ans_2_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_163 = _ans_2_leadingZeros_T_93[27] ? 6'h1b : _ans_2_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_164 = _ans_2_leadingZeros_T_93[26] ? 6'h1a : _ans_2_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_165 = _ans_2_leadingZeros_T_93[25] ? 6'h19 : _ans_2_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_166 = _ans_2_leadingZeros_T_93[24] ? 6'h18 : _ans_2_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_167 = _ans_2_leadingZeros_T_93[23] ? 6'h17 : _ans_2_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_168 = _ans_2_leadingZeros_T_93[22] ? 6'h16 : _ans_2_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_169 = _ans_2_leadingZeros_T_93[21] ? 6'h15 : _ans_2_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_170 = _ans_2_leadingZeros_T_93[20] ? 6'h14 : _ans_2_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_171 = _ans_2_leadingZeros_T_93[19] ? 6'h13 : _ans_2_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_172 = _ans_2_leadingZeros_T_93[18] ? 6'h12 : _ans_2_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_173 = _ans_2_leadingZeros_T_93[17] ? 6'h11 : _ans_2_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_174 = _ans_2_leadingZeros_T_93[16] ? 6'h10 : _ans_2_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_175 = _ans_2_leadingZeros_T_93[15] ? 6'hf : _ans_2_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_176 = _ans_2_leadingZeros_T_93[14] ? 6'he : _ans_2_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_177 = _ans_2_leadingZeros_T_93[13] ? 6'hd : _ans_2_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_178 = _ans_2_leadingZeros_T_93[12] ? 6'hc : _ans_2_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_179 = _ans_2_leadingZeros_T_93[11] ? 6'hb : _ans_2_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_180 = _ans_2_leadingZeros_T_93[10] ? 6'ha : _ans_2_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_181 = _ans_2_leadingZeros_T_93[9] ? 6'h9 : _ans_2_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_182 = _ans_2_leadingZeros_T_93[8] ? 6'h8 : _ans_2_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_183 = _ans_2_leadingZeros_T_93[7] ? 6'h7 : _ans_2_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_184 = _ans_2_leadingZeros_T_93[6] ? 6'h6 : _ans_2_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_185 = _ans_2_leadingZeros_T_93[5] ? 6'h5 : _ans_2_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_186 = _ans_2_leadingZeros_T_93[4] ? 6'h4 : _ans_2_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_187 = _ans_2_leadingZeros_T_93[3] ? 6'h3 : _ans_2_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_188 = _ans_2_leadingZeros_T_93[2] ? 6'h2 : _ans_2_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_189 = _ans_2_leadingZeros_T_93[1] ? 6'h1 : _ans_2_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_2_leadingZeros = _ans_2_leadingZeros_T_93[0] ? 6'h0 : _ans_2_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_expRaw_T_1 = 6'h1f - ans_2_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_2_expRaw = ans_2_isZero ? 6'h0 : _ans_2_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_2_shiftAmt_T_2 = ans_2_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_2_shiftAmt = ans_2_expRaw > 6'h3 ? _ans_2_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_2_mantissaRaw_T = ans_2_absClipped >> ans_2_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_2_mantissaRaw = _ans_2_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_2_mantissa = ans_2_expRaw >= 6'h3 ? ans_2_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_2_expAdjusted = ans_2_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_2_exp_T_4 = ans_2_expAdjusted > 7'hf ? 4'hf : ans_2_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_2_exp = ans_2_isZero ? 4'h0 : _ans_2_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_2_fp8 = {ans_2_clippedX[31],ans_2_exp,ans_2_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_3 = {24'h0,linear_bias_3}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_3 = tempSum_3 + biasExtended_3; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_3_sign = sum32_3[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_3_absX_T = ~sum32_3; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_3_absX_T_2 = _ans_3_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_3_absX = ans_3_sign ? _ans_3_absX_T_2 : sum32_3; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_3_shiftedX_T_1 = _GEN_10432 - ans_3_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_3_shiftedX_T_3 = ans_3_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_3_shiftedX = ans_3_sign ? _ans_3_shiftedX_T_1 : _ans_3_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_3_scaledX_T_1 = ans_3_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_3_scaledX = _ans_3_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_3_clippedX_T_2 = ans_3_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_3_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_3_clippedX = ans_3_scaledX > 49'h1c0 ? 49'h1c0 : _ans_3_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_3_absClipped_T_1 = ~ans_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_3_absClipped_T_3 = _ans_3_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_3_absClipped = ans_3_clippedX[31] ? _ans_3_absClipped_T_3 : ans_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_3_isZero = ans_3_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10467 = {{16'd0}, ans_3_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_4 = _GEN_10467 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_6 = {ans_3_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_8 = _ans_3_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_9 = _ans_3_leadingZeros_T_4 | _ans_3_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10468 = {{8'd0}, _ans_3_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_14 = _GEN_10468 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_16 = {_ans_3_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_18 = _ans_3_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_19 = _ans_3_leadingZeros_T_14 | _ans_3_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10469 = {{4'd0}, _ans_3_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_24 = _GEN_10469 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_26 = {_ans_3_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_28 = _ans_3_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_29 = _ans_3_leadingZeros_T_24 | _ans_3_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10470 = {{2'd0}, _ans_3_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_34 = _GEN_10470 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_36 = {_ans_3_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_38 = _ans_3_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_39 = _ans_3_leadingZeros_T_34 | _ans_3_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10471 = {{1'd0}, _ans_3_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_44 = _GEN_10471 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_46 = {_ans_3_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_48 = _ans_3_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_3_leadingZeros_T_49 = _ans_3_leadingZeros_T_44 | _ans_3_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10472 = {{8'd0}, ans_3_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_55 = _GEN_10472 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_57 = {ans_3_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_59 = _ans_3_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_60 = _ans_3_leadingZeros_T_55 | _ans_3_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10473 = {{4'd0}, _ans_3_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_65 = _GEN_10473 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_67 = {_ans_3_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_69 = _ans_3_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_70 = _ans_3_leadingZeros_T_65 | _ans_3_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10474 = {{2'd0}, _ans_3_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_75 = _GEN_10474 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_77 = {_ans_3_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_79 = _ans_3_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_80 = _ans_3_leadingZeros_T_75 | _ans_3_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10475 = {{1'd0}, _ans_3_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_85 = _GEN_10475 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_87 = {_ans_3_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_89 = _ans_3_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_3_leadingZeros_T_90 = _ans_3_leadingZeros_T_85 | _ans_3_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_3_leadingZeros_T_93 = {_ans_3_leadingZeros_T_49,_ans_3_leadingZeros_T_90,ans_3_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_3_leadingZeros_T_143 = _ans_3_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_144 = _ans_3_leadingZeros_T_93[46] ? 6'h2e : _ans_3_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_145 = _ans_3_leadingZeros_T_93[45] ? 6'h2d : _ans_3_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_146 = _ans_3_leadingZeros_T_93[44] ? 6'h2c : _ans_3_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_147 = _ans_3_leadingZeros_T_93[43] ? 6'h2b : _ans_3_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_148 = _ans_3_leadingZeros_T_93[42] ? 6'h2a : _ans_3_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_149 = _ans_3_leadingZeros_T_93[41] ? 6'h29 : _ans_3_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_150 = _ans_3_leadingZeros_T_93[40] ? 6'h28 : _ans_3_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_151 = _ans_3_leadingZeros_T_93[39] ? 6'h27 : _ans_3_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_152 = _ans_3_leadingZeros_T_93[38] ? 6'h26 : _ans_3_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_153 = _ans_3_leadingZeros_T_93[37] ? 6'h25 : _ans_3_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_154 = _ans_3_leadingZeros_T_93[36] ? 6'h24 : _ans_3_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_155 = _ans_3_leadingZeros_T_93[35] ? 6'h23 : _ans_3_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_156 = _ans_3_leadingZeros_T_93[34] ? 6'h22 : _ans_3_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_157 = _ans_3_leadingZeros_T_93[33] ? 6'h21 : _ans_3_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_158 = _ans_3_leadingZeros_T_93[32] ? 6'h20 : _ans_3_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_159 = _ans_3_leadingZeros_T_93[31] ? 6'h1f : _ans_3_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_160 = _ans_3_leadingZeros_T_93[30] ? 6'h1e : _ans_3_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_161 = _ans_3_leadingZeros_T_93[29] ? 6'h1d : _ans_3_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_162 = _ans_3_leadingZeros_T_93[28] ? 6'h1c : _ans_3_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_163 = _ans_3_leadingZeros_T_93[27] ? 6'h1b : _ans_3_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_164 = _ans_3_leadingZeros_T_93[26] ? 6'h1a : _ans_3_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_165 = _ans_3_leadingZeros_T_93[25] ? 6'h19 : _ans_3_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_166 = _ans_3_leadingZeros_T_93[24] ? 6'h18 : _ans_3_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_167 = _ans_3_leadingZeros_T_93[23] ? 6'h17 : _ans_3_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_168 = _ans_3_leadingZeros_T_93[22] ? 6'h16 : _ans_3_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_169 = _ans_3_leadingZeros_T_93[21] ? 6'h15 : _ans_3_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_170 = _ans_3_leadingZeros_T_93[20] ? 6'h14 : _ans_3_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_171 = _ans_3_leadingZeros_T_93[19] ? 6'h13 : _ans_3_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_172 = _ans_3_leadingZeros_T_93[18] ? 6'h12 : _ans_3_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_173 = _ans_3_leadingZeros_T_93[17] ? 6'h11 : _ans_3_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_174 = _ans_3_leadingZeros_T_93[16] ? 6'h10 : _ans_3_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_175 = _ans_3_leadingZeros_T_93[15] ? 6'hf : _ans_3_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_176 = _ans_3_leadingZeros_T_93[14] ? 6'he : _ans_3_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_177 = _ans_3_leadingZeros_T_93[13] ? 6'hd : _ans_3_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_178 = _ans_3_leadingZeros_T_93[12] ? 6'hc : _ans_3_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_179 = _ans_3_leadingZeros_T_93[11] ? 6'hb : _ans_3_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_180 = _ans_3_leadingZeros_T_93[10] ? 6'ha : _ans_3_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_181 = _ans_3_leadingZeros_T_93[9] ? 6'h9 : _ans_3_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_182 = _ans_3_leadingZeros_T_93[8] ? 6'h8 : _ans_3_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_183 = _ans_3_leadingZeros_T_93[7] ? 6'h7 : _ans_3_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_184 = _ans_3_leadingZeros_T_93[6] ? 6'h6 : _ans_3_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_185 = _ans_3_leadingZeros_T_93[5] ? 6'h5 : _ans_3_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_186 = _ans_3_leadingZeros_T_93[4] ? 6'h4 : _ans_3_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_187 = _ans_3_leadingZeros_T_93[3] ? 6'h3 : _ans_3_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_188 = _ans_3_leadingZeros_T_93[2] ? 6'h2 : _ans_3_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_189 = _ans_3_leadingZeros_T_93[1] ? 6'h1 : _ans_3_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_3_leadingZeros = _ans_3_leadingZeros_T_93[0] ? 6'h0 : _ans_3_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_expRaw_T_1 = 6'h1f - ans_3_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_3_expRaw = ans_3_isZero ? 6'h0 : _ans_3_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_3_shiftAmt_T_2 = ans_3_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_3_shiftAmt = ans_3_expRaw > 6'h3 ? _ans_3_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_3_mantissaRaw_T = ans_3_absClipped >> ans_3_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_3_mantissaRaw = _ans_3_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_3_mantissa = ans_3_expRaw >= 6'h3 ? ans_3_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_3_expAdjusted = ans_3_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_3_exp_T_4 = ans_3_expAdjusted > 7'hf ? 4'hf : ans_3_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_3_exp = ans_3_isZero ? 4'h0 : _ans_3_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_3_fp8 = {ans_3_clippedX[31],ans_3_exp,ans_3_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_4 = {24'h0,linear_bias_4}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_4 = tempSum_4 + biasExtended_4; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_4_sign = sum32_4[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_4_absX_T = ~sum32_4; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_4_absX_T_2 = _ans_4_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_4_absX = ans_4_sign ? _ans_4_absX_T_2 : sum32_4; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_4_shiftedX_T_1 = _GEN_10432 - ans_4_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_4_shiftedX_T_3 = ans_4_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_4_shiftedX = ans_4_sign ? _ans_4_shiftedX_T_1 : _ans_4_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_4_scaledX_T_1 = ans_4_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_4_scaledX = _ans_4_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_4_clippedX_T_2 = ans_4_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_4_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_4_clippedX = ans_4_scaledX > 49'h1c0 ? 49'h1c0 : _ans_4_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_4_absClipped_T_1 = ~ans_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_4_absClipped_T_3 = _ans_4_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_4_absClipped = ans_4_clippedX[31] ? _ans_4_absClipped_T_3 : ans_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_4_isZero = ans_4_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10478 = {{16'd0}, ans_4_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_4 = _GEN_10478 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_6 = {ans_4_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_8 = _ans_4_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_9 = _ans_4_leadingZeros_T_4 | _ans_4_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10479 = {{8'd0}, _ans_4_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_14 = _GEN_10479 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_16 = {_ans_4_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_18 = _ans_4_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_19 = _ans_4_leadingZeros_T_14 | _ans_4_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10480 = {{4'd0}, _ans_4_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_24 = _GEN_10480 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_26 = {_ans_4_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_28 = _ans_4_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_29 = _ans_4_leadingZeros_T_24 | _ans_4_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10481 = {{2'd0}, _ans_4_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_34 = _GEN_10481 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_36 = {_ans_4_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_38 = _ans_4_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_39 = _ans_4_leadingZeros_T_34 | _ans_4_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10482 = {{1'd0}, _ans_4_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_44 = _GEN_10482 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_46 = {_ans_4_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_48 = _ans_4_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_4_leadingZeros_T_49 = _ans_4_leadingZeros_T_44 | _ans_4_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10483 = {{8'd0}, ans_4_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_55 = _GEN_10483 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_57 = {ans_4_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_59 = _ans_4_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_60 = _ans_4_leadingZeros_T_55 | _ans_4_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10484 = {{4'd0}, _ans_4_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_65 = _GEN_10484 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_67 = {_ans_4_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_69 = _ans_4_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_70 = _ans_4_leadingZeros_T_65 | _ans_4_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10485 = {{2'd0}, _ans_4_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_75 = _GEN_10485 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_77 = {_ans_4_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_79 = _ans_4_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_80 = _ans_4_leadingZeros_T_75 | _ans_4_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10486 = {{1'd0}, _ans_4_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_85 = _GEN_10486 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_87 = {_ans_4_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_89 = _ans_4_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_4_leadingZeros_T_90 = _ans_4_leadingZeros_T_85 | _ans_4_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_4_leadingZeros_T_93 = {_ans_4_leadingZeros_T_49,_ans_4_leadingZeros_T_90,ans_4_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_4_leadingZeros_T_143 = _ans_4_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_144 = _ans_4_leadingZeros_T_93[46] ? 6'h2e : _ans_4_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_145 = _ans_4_leadingZeros_T_93[45] ? 6'h2d : _ans_4_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_146 = _ans_4_leadingZeros_T_93[44] ? 6'h2c : _ans_4_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_147 = _ans_4_leadingZeros_T_93[43] ? 6'h2b : _ans_4_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_148 = _ans_4_leadingZeros_T_93[42] ? 6'h2a : _ans_4_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_149 = _ans_4_leadingZeros_T_93[41] ? 6'h29 : _ans_4_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_150 = _ans_4_leadingZeros_T_93[40] ? 6'h28 : _ans_4_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_151 = _ans_4_leadingZeros_T_93[39] ? 6'h27 : _ans_4_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_152 = _ans_4_leadingZeros_T_93[38] ? 6'h26 : _ans_4_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_153 = _ans_4_leadingZeros_T_93[37] ? 6'h25 : _ans_4_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_154 = _ans_4_leadingZeros_T_93[36] ? 6'h24 : _ans_4_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_155 = _ans_4_leadingZeros_T_93[35] ? 6'h23 : _ans_4_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_156 = _ans_4_leadingZeros_T_93[34] ? 6'h22 : _ans_4_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_157 = _ans_4_leadingZeros_T_93[33] ? 6'h21 : _ans_4_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_158 = _ans_4_leadingZeros_T_93[32] ? 6'h20 : _ans_4_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_159 = _ans_4_leadingZeros_T_93[31] ? 6'h1f : _ans_4_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_160 = _ans_4_leadingZeros_T_93[30] ? 6'h1e : _ans_4_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_161 = _ans_4_leadingZeros_T_93[29] ? 6'h1d : _ans_4_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_162 = _ans_4_leadingZeros_T_93[28] ? 6'h1c : _ans_4_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_163 = _ans_4_leadingZeros_T_93[27] ? 6'h1b : _ans_4_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_164 = _ans_4_leadingZeros_T_93[26] ? 6'h1a : _ans_4_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_165 = _ans_4_leadingZeros_T_93[25] ? 6'h19 : _ans_4_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_166 = _ans_4_leadingZeros_T_93[24] ? 6'h18 : _ans_4_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_167 = _ans_4_leadingZeros_T_93[23] ? 6'h17 : _ans_4_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_168 = _ans_4_leadingZeros_T_93[22] ? 6'h16 : _ans_4_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_169 = _ans_4_leadingZeros_T_93[21] ? 6'h15 : _ans_4_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_170 = _ans_4_leadingZeros_T_93[20] ? 6'h14 : _ans_4_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_171 = _ans_4_leadingZeros_T_93[19] ? 6'h13 : _ans_4_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_172 = _ans_4_leadingZeros_T_93[18] ? 6'h12 : _ans_4_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_173 = _ans_4_leadingZeros_T_93[17] ? 6'h11 : _ans_4_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_174 = _ans_4_leadingZeros_T_93[16] ? 6'h10 : _ans_4_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_175 = _ans_4_leadingZeros_T_93[15] ? 6'hf : _ans_4_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_176 = _ans_4_leadingZeros_T_93[14] ? 6'he : _ans_4_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_177 = _ans_4_leadingZeros_T_93[13] ? 6'hd : _ans_4_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_178 = _ans_4_leadingZeros_T_93[12] ? 6'hc : _ans_4_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_179 = _ans_4_leadingZeros_T_93[11] ? 6'hb : _ans_4_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_180 = _ans_4_leadingZeros_T_93[10] ? 6'ha : _ans_4_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_181 = _ans_4_leadingZeros_T_93[9] ? 6'h9 : _ans_4_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_182 = _ans_4_leadingZeros_T_93[8] ? 6'h8 : _ans_4_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_183 = _ans_4_leadingZeros_T_93[7] ? 6'h7 : _ans_4_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_184 = _ans_4_leadingZeros_T_93[6] ? 6'h6 : _ans_4_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_185 = _ans_4_leadingZeros_T_93[5] ? 6'h5 : _ans_4_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_186 = _ans_4_leadingZeros_T_93[4] ? 6'h4 : _ans_4_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_187 = _ans_4_leadingZeros_T_93[3] ? 6'h3 : _ans_4_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_188 = _ans_4_leadingZeros_T_93[2] ? 6'h2 : _ans_4_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_189 = _ans_4_leadingZeros_T_93[1] ? 6'h1 : _ans_4_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_4_leadingZeros = _ans_4_leadingZeros_T_93[0] ? 6'h0 : _ans_4_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_expRaw_T_1 = 6'h1f - ans_4_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_4_expRaw = ans_4_isZero ? 6'h0 : _ans_4_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_4_shiftAmt_T_2 = ans_4_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_4_shiftAmt = ans_4_expRaw > 6'h3 ? _ans_4_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_4_mantissaRaw_T = ans_4_absClipped >> ans_4_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_4_mantissaRaw = _ans_4_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_4_mantissa = ans_4_expRaw >= 6'h3 ? ans_4_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_4_expAdjusted = ans_4_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_4_exp_T_4 = ans_4_expAdjusted > 7'hf ? 4'hf : ans_4_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_4_exp = ans_4_isZero ? 4'h0 : _ans_4_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_4_fp8 = {ans_4_clippedX[31],ans_4_exp,ans_4_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_5 = {24'h0,linear_bias_5}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_5 = tempSum_5 + biasExtended_5; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_5_sign = sum32_5[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_5_absX_T = ~sum32_5; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_5_absX_T_2 = _ans_5_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_5_absX = ans_5_sign ? _ans_5_absX_T_2 : sum32_5; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_5_shiftedX_T_1 = _GEN_10432 - ans_5_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_5_shiftedX_T_3 = ans_5_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_5_shiftedX = ans_5_sign ? _ans_5_shiftedX_T_1 : _ans_5_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_5_scaledX_T_1 = ans_5_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_5_scaledX = _ans_5_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_5_clippedX_T_2 = ans_5_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_5_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_5_clippedX = ans_5_scaledX > 49'h1c0 ? 49'h1c0 : _ans_5_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_5_absClipped_T_1 = ~ans_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_5_absClipped_T_3 = _ans_5_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_5_absClipped = ans_5_clippedX[31] ? _ans_5_absClipped_T_3 : ans_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_5_isZero = ans_5_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10489 = {{16'd0}, ans_5_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_4 = _GEN_10489 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_6 = {ans_5_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_8 = _ans_5_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_9 = _ans_5_leadingZeros_T_4 | _ans_5_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10490 = {{8'd0}, _ans_5_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_14 = _GEN_10490 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_16 = {_ans_5_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_18 = _ans_5_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_19 = _ans_5_leadingZeros_T_14 | _ans_5_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10491 = {{4'd0}, _ans_5_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_24 = _GEN_10491 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_26 = {_ans_5_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_28 = _ans_5_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_29 = _ans_5_leadingZeros_T_24 | _ans_5_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10492 = {{2'd0}, _ans_5_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_34 = _GEN_10492 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_36 = {_ans_5_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_38 = _ans_5_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_39 = _ans_5_leadingZeros_T_34 | _ans_5_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10493 = {{1'd0}, _ans_5_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_44 = _GEN_10493 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_46 = {_ans_5_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_48 = _ans_5_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_5_leadingZeros_T_49 = _ans_5_leadingZeros_T_44 | _ans_5_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10494 = {{8'd0}, ans_5_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_55 = _GEN_10494 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_57 = {ans_5_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_59 = _ans_5_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_60 = _ans_5_leadingZeros_T_55 | _ans_5_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10495 = {{4'd0}, _ans_5_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_65 = _GEN_10495 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_67 = {_ans_5_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_69 = _ans_5_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_70 = _ans_5_leadingZeros_T_65 | _ans_5_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10496 = {{2'd0}, _ans_5_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_75 = _GEN_10496 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_77 = {_ans_5_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_79 = _ans_5_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_80 = _ans_5_leadingZeros_T_75 | _ans_5_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10497 = {{1'd0}, _ans_5_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_85 = _GEN_10497 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_87 = {_ans_5_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_89 = _ans_5_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_5_leadingZeros_T_90 = _ans_5_leadingZeros_T_85 | _ans_5_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_5_leadingZeros_T_93 = {_ans_5_leadingZeros_T_49,_ans_5_leadingZeros_T_90,ans_5_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_5_leadingZeros_T_143 = _ans_5_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_144 = _ans_5_leadingZeros_T_93[46] ? 6'h2e : _ans_5_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_145 = _ans_5_leadingZeros_T_93[45] ? 6'h2d : _ans_5_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_146 = _ans_5_leadingZeros_T_93[44] ? 6'h2c : _ans_5_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_147 = _ans_5_leadingZeros_T_93[43] ? 6'h2b : _ans_5_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_148 = _ans_5_leadingZeros_T_93[42] ? 6'h2a : _ans_5_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_149 = _ans_5_leadingZeros_T_93[41] ? 6'h29 : _ans_5_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_150 = _ans_5_leadingZeros_T_93[40] ? 6'h28 : _ans_5_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_151 = _ans_5_leadingZeros_T_93[39] ? 6'h27 : _ans_5_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_152 = _ans_5_leadingZeros_T_93[38] ? 6'h26 : _ans_5_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_153 = _ans_5_leadingZeros_T_93[37] ? 6'h25 : _ans_5_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_154 = _ans_5_leadingZeros_T_93[36] ? 6'h24 : _ans_5_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_155 = _ans_5_leadingZeros_T_93[35] ? 6'h23 : _ans_5_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_156 = _ans_5_leadingZeros_T_93[34] ? 6'h22 : _ans_5_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_157 = _ans_5_leadingZeros_T_93[33] ? 6'h21 : _ans_5_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_158 = _ans_5_leadingZeros_T_93[32] ? 6'h20 : _ans_5_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_159 = _ans_5_leadingZeros_T_93[31] ? 6'h1f : _ans_5_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_160 = _ans_5_leadingZeros_T_93[30] ? 6'h1e : _ans_5_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_161 = _ans_5_leadingZeros_T_93[29] ? 6'h1d : _ans_5_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_162 = _ans_5_leadingZeros_T_93[28] ? 6'h1c : _ans_5_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_163 = _ans_5_leadingZeros_T_93[27] ? 6'h1b : _ans_5_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_164 = _ans_5_leadingZeros_T_93[26] ? 6'h1a : _ans_5_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_165 = _ans_5_leadingZeros_T_93[25] ? 6'h19 : _ans_5_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_166 = _ans_5_leadingZeros_T_93[24] ? 6'h18 : _ans_5_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_167 = _ans_5_leadingZeros_T_93[23] ? 6'h17 : _ans_5_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_168 = _ans_5_leadingZeros_T_93[22] ? 6'h16 : _ans_5_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_169 = _ans_5_leadingZeros_T_93[21] ? 6'h15 : _ans_5_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_170 = _ans_5_leadingZeros_T_93[20] ? 6'h14 : _ans_5_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_171 = _ans_5_leadingZeros_T_93[19] ? 6'h13 : _ans_5_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_172 = _ans_5_leadingZeros_T_93[18] ? 6'h12 : _ans_5_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_173 = _ans_5_leadingZeros_T_93[17] ? 6'h11 : _ans_5_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_174 = _ans_5_leadingZeros_T_93[16] ? 6'h10 : _ans_5_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_175 = _ans_5_leadingZeros_T_93[15] ? 6'hf : _ans_5_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_176 = _ans_5_leadingZeros_T_93[14] ? 6'he : _ans_5_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_177 = _ans_5_leadingZeros_T_93[13] ? 6'hd : _ans_5_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_178 = _ans_5_leadingZeros_T_93[12] ? 6'hc : _ans_5_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_179 = _ans_5_leadingZeros_T_93[11] ? 6'hb : _ans_5_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_180 = _ans_5_leadingZeros_T_93[10] ? 6'ha : _ans_5_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_181 = _ans_5_leadingZeros_T_93[9] ? 6'h9 : _ans_5_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_182 = _ans_5_leadingZeros_T_93[8] ? 6'h8 : _ans_5_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_183 = _ans_5_leadingZeros_T_93[7] ? 6'h7 : _ans_5_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_184 = _ans_5_leadingZeros_T_93[6] ? 6'h6 : _ans_5_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_185 = _ans_5_leadingZeros_T_93[5] ? 6'h5 : _ans_5_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_186 = _ans_5_leadingZeros_T_93[4] ? 6'h4 : _ans_5_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_187 = _ans_5_leadingZeros_T_93[3] ? 6'h3 : _ans_5_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_188 = _ans_5_leadingZeros_T_93[2] ? 6'h2 : _ans_5_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_189 = _ans_5_leadingZeros_T_93[1] ? 6'h1 : _ans_5_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_5_leadingZeros = _ans_5_leadingZeros_T_93[0] ? 6'h0 : _ans_5_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_expRaw_T_1 = 6'h1f - ans_5_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_5_expRaw = ans_5_isZero ? 6'h0 : _ans_5_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_5_shiftAmt_T_2 = ans_5_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_5_shiftAmt = ans_5_expRaw > 6'h3 ? _ans_5_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_5_mantissaRaw_T = ans_5_absClipped >> ans_5_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_5_mantissaRaw = _ans_5_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_5_mantissa = ans_5_expRaw >= 6'h3 ? ans_5_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_5_expAdjusted = ans_5_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_5_exp_T_4 = ans_5_expAdjusted > 7'hf ? 4'hf : ans_5_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_5_exp = ans_5_isZero ? 4'h0 : _ans_5_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_5_fp8 = {ans_5_clippedX[31],ans_5_exp,ans_5_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_6 = {24'h0,linear_bias_6}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_6 = tempSum_6 + biasExtended_6; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_6_sign = sum32_6[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_6_absX_T = ~sum32_6; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_6_absX_T_2 = _ans_6_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_6_absX = ans_6_sign ? _ans_6_absX_T_2 : sum32_6; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_6_shiftedX_T_1 = _GEN_10432 - ans_6_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_6_shiftedX_T_3 = ans_6_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_6_shiftedX = ans_6_sign ? _ans_6_shiftedX_T_1 : _ans_6_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_6_scaledX_T_1 = ans_6_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_6_scaledX = _ans_6_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_6_clippedX_T_2 = ans_6_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_6_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_6_clippedX = ans_6_scaledX > 49'h1c0 ? 49'h1c0 : _ans_6_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_6_absClipped_T_1 = ~ans_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_6_absClipped_T_3 = _ans_6_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_6_absClipped = ans_6_clippedX[31] ? _ans_6_absClipped_T_3 : ans_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_6_isZero = ans_6_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10500 = {{16'd0}, ans_6_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_4 = _GEN_10500 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_6 = {ans_6_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_8 = _ans_6_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_9 = _ans_6_leadingZeros_T_4 | _ans_6_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10501 = {{8'd0}, _ans_6_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_14 = _GEN_10501 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_16 = {_ans_6_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_18 = _ans_6_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_19 = _ans_6_leadingZeros_T_14 | _ans_6_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10502 = {{4'd0}, _ans_6_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_24 = _GEN_10502 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_26 = {_ans_6_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_28 = _ans_6_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_29 = _ans_6_leadingZeros_T_24 | _ans_6_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10503 = {{2'd0}, _ans_6_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_34 = _GEN_10503 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_36 = {_ans_6_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_38 = _ans_6_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_39 = _ans_6_leadingZeros_T_34 | _ans_6_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10504 = {{1'd0}, _ans_6_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_44 = _GEN_10504 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_46 = {_ans_6_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_48 = _ans_6_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_6_leadingZeros_T_49 = _ans_6_leadingZeros_T_44 | _ans_6_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10505 = {{8'd0}, ans_6_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_55 = _GEN_10505 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_57 = {ans_6_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_59 = _ans_6_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_60 = _ans_6_leadingZeros_T_55 | _ans_6_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10506 = {{4'd0}, _ans_6_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_65 = _GEN_10506 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_67 = {_ans_6_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_69 = _ans_6_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_70 = _ans_6_leadingZeros_T_65 | _ans_6_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10507 = {{2'd0}, _ans_6_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_75 = _GEN_10507 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_77 = {_ans_6_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_79 = _ans_6_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_80 = _ans_6_leadingZeros_T_75 | _ans_6_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10508 = {{1'd0}, _ans_6_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_85 = _GEN_10508 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_87 = {_ans_6_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_89 = _ans_6_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_6_leadingZeros_T_90 = _ans_6_leadingZeros_T_85 | _ans_6_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_6_leadingZeros_T_93 = {_ans_6_leadingZeros_T_49,_ans_6_leadingZeros_T_90,ans_6_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_6_leadingZeros_T_143 = _ans_6_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_144 = _ans_6_leadingZeros_T_93[46] ? 6'h2e : _ans_6_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_145 = _ans_6_leadingZeros_T_93[45] ? 6'h2d : _ans_6_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_146 = _ans_6_leadingZeros_T_93[44] ? 6'h2c : _ans_6_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_147 = _ans_6_leadingZeros_T_93[43] ? 6'h2b : _ans_6_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_148 = _ans_6_leadingZeros_T_93[42] ? 6'h2a : _ans_6_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_149 = _ans_6_leadingZeros_T_93[41] ? 6'h29 : _ans_6_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_150 = _ans_6_leadingZeros_T_93[40] ? 6'h28 : _ans_6_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_151 = _ans_6_leadingZeros_T_93[39] ? 6'h27 : _ans_6_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_152 = _ans_6_leadingZeros_T_93[38] ? 6'h26 : _ans_6_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_153 = _ans_6_leadingZeros_T_93[37] ? 6'h25 : _ans_6_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_154 = _ans_6_leadingZeros_T_93[36] ? 6'h24 : _ans_6_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_155 = _ans_6_leadingZeros_T_93[35] ? 6'h23 : _ans_6_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_156 = _ans_6_leadingZeros_T_93[34] ? 6'h22 : _ans_6_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_157 = _ans_6_leadingZeros_T_93[33] ? 6'h21 : _ans_6_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_158 = _ans_6_leadingZeros_T_93[32] ? 6'h20 : _ans_6_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_159 = _ans_6_leadingZeros_T_93[31] ? 6'h1f : _ans_6_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_160 = _ans_6_leadingZeros_T_93[30] ? 6'h1e : _ans_6_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_161 = _ans_6_leadingZeros_T_93[29] ? 6'h1d : _ans_6_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_162 = _ans_6_leadingZeros_T_93[28] ? 6'h1c : _ans_6_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_163 = _ans_6_leadingZeros_T_93[27] ? 6'h1b : _ans_6_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_164 = _ans_6_leadingZeros_T_93[26] ? 6'h1a : _ans_6_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_165 = _ans_6_leadingZeros_T_93[25] ? 6'h19 : _ans_6_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_166 = _ans_6_leadingZeros_T_93[24] ? 6'h18 : _ans_6_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_167 = _ans_6_leadingZeros_T_93[23] ? 6'h17 : _ans_6_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_168 = _ans_6_leadingZeros_T_93[22] ? 6'h16 : _ans_6_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_169 = _ans_6_leadingZeros_T_93[21] ? 6'h15 : _ans_6_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_170 = _ans_6_leadingZeros_T_93[20] ? 6'h14 : _ans_6_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_171 = _ans_6_leadingZeros_T_93[19] ? 6'h13 : _ans_6_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_172 = _ans_6_leadingZeros_T_93[18] ? 6'h12 : _ans_6_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_173 = _ans_6_leadingZeros_T_93[17] ? 6'h11 : _ans_6_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_174 = _ans_6_leadingZeros_T_93[16] ? 6'h10 : _ans_6_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_175 = _ans_6_leadingZeros_T_93[15] ? 6'hf : _ans_6_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_176 = _ans_6_leadingZeros_T_93[14] ? 6'he : _ans_6_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_177 = _ans_6_leadingZeros_T_93[13] ? 6'hd : _ans_6_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_178 = _ans_6_leadingZeros_T_93[12] ? 6'hc : _ans_6_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_179 = _ans_6_leadingZeros_T_93[11] ? 6'hb : _ans_6_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_180 = _ans_6_leadingZeros_T_93[10] ? 6'ha : _ans_6_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_181 = _ans_6_leadingZeros_T_93[9] ? 6'h9 : _ans_6_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_182 = _ans_6_leadingZeros_T_93[8] ? 6'h8 : _ans_6_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_183 = _ans_6_leadingZeros_T_93[7] ? 6'h7 : _ans_6_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_184 = _ans_6_leadingZeros_T_93[6] ? 6'h6 : _ans_6_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_185 = _ans_6_leadingZeros_T_93[5] ? 6'h5 : _ans_6_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_186 = _ans_6_leadingZeros_T_93[4] ? 6'h4 : _ans_6_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_187 = _ans_6_leadingZeros_T_93[3] ? 6'h3 : _ans_6_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_188 = _ans_6_leadingZeros_T_93[2] ? 6'h2 : _ans_6_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_189 = _ans_6_leadingZeros_T_93[1] ? 6'h1 : _ans_6_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_6_leadingZeros = _ans_6_leadingZeros_T_93[0] ? 6'h0 : _ans_6_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_expRaw_T_1 = 6'h1f - ans_6_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_6_expRaw = ans_6_isZero ? 6'h0 : _ans_6_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_6_shiftAmt_T_2 = ans_6_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_6_shiftAmt = ans_6_expRaw > 6'h3 ? _ans_6_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_6_mantissaRaw_T = ans_6_absClipped >> ans_6_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_6_mantissaRaw = _ans_6_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_6_mantissa = ans_6_expRaw >= 6'h3 ? ans_6_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_6_expAdjusted = ans_6_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_6_exp_T_4 = ans_6_expAdjusted > 7'hf ? 4'hf : ans_6_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_6_exp = ans_6_isZero ? 4'h0 : _ans_6_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_6_fp8 = {ans_6_clippedX[31],ans_6_exp,ans_6_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_7 = {24'h0,linear_bias_7}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_7 = tempSum_7 + biasExtended_7; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_7_sign = sum32_7[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_7_absX_T = ~sum32_7; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_7_absX_T_2 = _ans_7_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_7_absX = ans_7_sign ? _ans_7_absX_T_2 : sum32_7; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_7_shiftedX_T_1 = _GEN_10432 - ans_7_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_7_shiftedX_T_3 = ans_7_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_7_shiftedX = ans_7_sign ? _ans_7_shiftedX_T_1 : _ans_7_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_7_scaledX_T_1 = ans_7_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_7_scaledX = _ans_7_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_7_clippedX_T_2 = ans_7_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_7_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_7_clippedX = ans_7_scaledX > 49'h1c0 ? 49'h1c0 : _ans_7_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_7_absClipped_T_1 = ~ans_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_7_absClipped_T_3 = _ans_7_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_7_absClipped = ans_7_clippedX[31] ? _ans_7_absClipped_T_3 : ans_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_7_isZero = ans_7_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10511 = {{16'd0}, ans_7_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_4 = _GEN_10511 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_6 = {ans_7_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_8 = _ans_7_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_9 = _ans_7_leadingZeros_T_4 | _ans_7_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10512 = {{8'd0}, _ans_7_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_14 = _GEN_10512 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_16 = {_ans_7_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_18 = _ans_7_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_19 = _ans_7_leadingZeros_T_14 | _ans_7_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10513 = {{4'd0}, _ans_7_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_24 = _GEN_10513 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_26 = {_ans_7_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_28 = _ans_7_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_29 = _ans_7_leadingZeros_T_24 | _ans_7_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10514 = {{2'd0}, _ans_7_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_34 = _GEN_10514 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_36 = {_ans_7_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_38 = _ans_7_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_39 = _ans_7_leadingZeros_T_34 | _ans_7_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10515 = {{1'd0}, _ans_7_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_44 = _GEN_10515 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_46 = {_ans_7_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_48 = _ans_7_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_7_leadingZeros_T_49 = _ans_7_leadingZeros_T_44 | _ans_7_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10516 = {{8'd0}, ans_7_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_55 = _GEN_10516 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_57 = {ans_7_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_59 = _ans_7_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_60 = _ans_7_leadingZeros_T_55 | _ans_7_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10517 = {{4'd0}, _ans_7_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_65 = _GEN_10517 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_67 = {_ans_7_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_69 = _ans_7_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_70 = _ans_7_leadingZeros_T_65 | _ans_7_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10518 = {{2'd0}, _ans_7_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_75 = _GEN_10518 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_77 = {_ans_7_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_79 = _ans_7_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_80 = _ans_7_leadingZeros_T_75 | _ans_7_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10519 = {{1'd0}, _ans_7_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_85 = _GEN_10519 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_87 = {_ans_7_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_89 = _ans_7_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_7_leadingZeros_T_90 = _ans_7_leadingZeros_T_85 | _ans_7_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_7_leadingZeros_T_93 = {_ans_7_leadingZeros_T_49,_ans_7_leadingZeros_T_90,ans_7_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_7_leadingZeros_T_143 = _ans_7_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_144 = _ans_7_leadingZeros_T_93[46] ? 6'h2e : _ans_7_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_145 = _ans_7_leadingZeros_T_93[45] ? 6'h2d : _ans_7_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_146 = _ans_7_leadingZeros_T_93[44] ? 6'h2c : _ans_7_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_147 = _ans_7_leadingZeros_T_93[43] ? 6'h2b : _ans_7_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_148 = _ans_7_leadingZeros_T_93[42] ? 6'h2a : _ans_7_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_149 = _ans_7_leadingZeros_T_93[41] ? 6'h29 : _ans_7_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_150 = _ans_7_leadingZeros_T_93[40] ? 6'h28 : _ans_7_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_151 = _ans_7_leadingZeros_T_93[39] ? 6'h27 : _ans_7_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_152 = _ans_7_leadingZeros_T_93[38] ? 6'h26 : _ans_7_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_153 = _ans_7_leadingZeros_T_93[37] ? 6'h25 : _ans_7_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_154 = _ans_7_leadingZeros_T_93[36] ? 6'h24 : _ans_7_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_155 = _ans_7_leadingZeros_T_93[35] ? 6'h23 : _ans_7_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_156 = _ans_7_leadingZeros_T_93[34] ? 6'h22 : _ans_7_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_157 = _ans_7_leadingZeros_T_93[33] ? 6'h21 : _ans_7_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_158 = _ans_7_leadingZeros_T_93[32] ? 6'h20 : _ans_7_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_159 = _ans_7_leadingZeros_T_93[31] ? 6'h1f : _ans_7_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_160 = _ans_7_leadingZeros_T_93[30] ? 6'h1e : _ans_7_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_161 = _ans_7_leadingZeros_T_93[29] ? 6'h1d : _ans_7_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_162 = _ans_7_leadingZeros_T_93[28] ? 6'h1c : _ans_7_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_163 = _ans_7_leadingZeros_T_93[27] ? 6'h1b : _ans_7_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_164 = _ans_7_leadingZeros_T_93[26] ? 6'h1a : _ans_7_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_165 = _ans_7_leadingZeros_T_93[25] ? 6'h19 : _ans_7_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_166 = _ans_7_leadingZeros_T_93[24] ? 6'h18 : _ans_7_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_167 = _ans_7_leadingZeros_T_93[23] ? 6'h17 : _ans_7_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_168 = _ans_7_leadingZeros_T_93[22] ? 6'h16 : _ans_7_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_169 = _ans_7_leadingZeros_T_93[21] ? 6'h15 : _ans_7_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_170 = _ans_7_leadingZeros_T_93[20] ? 6'h14 : _ans_7_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_171 = _ans_7_leadingZeros_T_93[19] ? 6'h13 : _ans_7_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_172 = _ans_7_leadingZeros_T_93[18] ? 6'h12 : _ans_7_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_173 = _ans_7_leadingZeros_T_93[17] ? 6'h11 : _ans_7_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_174 = _ans_7_leadingZeros_T_93[16] ? 6'h10 : _ans_7_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_175 = _ans_7_leadingZeros_T_93[15] ? 6'hf : _ans_7_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_176 = _ans_7_leadingZeros_T_93[14] ? 6'he : _ans_7_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_177 = _ans_7_leadingZeros_T_93[13] ? 6'hd : _ans_7_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_178 = _ans_7_leadingZeros_T_93[12] ? 6'hc : _ans_7_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_179 = _ans_7_leadingZeros_T_93[11] ? 6'hb : _ans_7_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_180 = _ans_7_leadingZeros_T_93[10] ? 6'ha : _ans_7_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_181 = _ans_7_leadingZeros_T_93[9] ? 6'h9 : _ans_7_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_182 = _ans_7_leadingZeros_T_93[8] ? 6'h8 : _ans_7_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_183 = _ans_7_leadingZeros_T_93[7] ? 6'h7 : _ans_7_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_184 = _ans_7_leadingZeros_T_93[6] ? 6'h6 : _ans_7_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_185 = _ans_7_leadingZeros_T_93[5] ? 6'h5 : _ans_7_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_186 = _ans_7_leadingZeros_T_93[4] ? 6'h4 : _ans_7_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_187 = _ans_7_leadingZeros_T_93[3] ? 6'h3 : _ans_7_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_188 = _ans_7_leadingZeros_T_93[2] ? 6'h2 : _ans_7_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_189 = _ans_7_leadingZeros_T_93[1] ? 6'h1 : _ans_7_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_7_leadingZeros = _ans_7_leadingZeros_T_93[0] ? 6'h0 : _ans_7_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_expRaw_T_1 = 6'h1f - ans_7_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_7_expRaw = ans_7_isZero ? 6'h0 : _ans_7_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_7_shiftAmt_T_2 = ans_7_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_7_shiftAmt = ans_7_expRaw > 6'h3 ? _ans_7_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_7_mantissaRaw_T = ans_7_absClipped >> ans_7_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_7_mantissaRaw = _ans_7_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_7_mantissa = ans_7_expRaw >= 6'h3 ? ans_7_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_7_expAdjusted = ans_7_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_7_exp_T_4 = ans_7_expAdjusted > 7'hf ? 4'hf : ans_7_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_7_exp = ans_7_isZero ? 4'h0 : _ans_7_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_7_fp8 = {ans_7_clippedX[31],ans_7_exp,ans_7_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_8 = {24'h0,linear_bias_8}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_8 = tempSum_8 + biasExtended_8; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_8_sign = sum32_8[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_8_absX_T = ~sum32_8; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_8_absX_T_2 = _ans_8_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_8_absX = ans_8_sign ? _ans_8_absX_T_2 : sum32_8; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_8_shiftedX_T_1 = _GEN_10432 - ans_8_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_8_shiftedX_T_3 = ans_8_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_8_shiftedX = ans_8_sign ? _ans_8_shiftedX_T_1 : _ans_8_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_8_scaledX_T_1 = ans_8_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_8_scaledX = _ans_8_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_8_clippedX_T_2 = ans_8_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_8_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_8_clippedX = ans_8_scaledX > 49'h1c0 ? 49'h1c0 : _ans_8_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_8_absClipped_T_1 = ~ans_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_8_absClipped_T_3 = _ans_8_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_8_absClipped = ans_8_clippedX[31] ? _ans_8_absClipped_T_3 : ans_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_8_isZero = ans_8_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10522 = {{16'd0}, ans_8_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_4 = _GEN_10522 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_6 = {ans_8_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_8 = _ans_8_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_9 = _ans_8_leadingZeros_T_4 | _ans_8_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10523 = {{8'd0}, _ans_8_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_14 = _GEN_10523 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_16 = {_ans_8_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_18 = _ans_8_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_19 = _ans_8_leadingZeros_T_14 | _ans_8_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10524 = {{4'd0}, _ans_8_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_24 = _GEN_10524 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_26 = {_ans_8_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_28 = _ans_8_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_29 = _ans_8_leadingZeros_T_24 | _ans_8_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10525 = {{2'd0}, _ans_8_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_34 = _GEN_10525 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_36 = {_ans_8_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_38 = _ans_8_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_39 = _ans_8_leadingZeros_T_34 | _ans_8_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10526 = {{1'd0}, _ans_8_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_44 = _GEN_10526 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_46 = {_ans_8_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_48 = _ans_8_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_8_leadingZeros_T_49 = _ans_8_leadingZeros_T_44 | _ans_8_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10527 = {{8'd0}, ans_8_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_55 = _GEN_10527 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_57 = {ans_8_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_59 = _ans_8_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_60 = _ans_8_leadingZeros_T_55 | _ans_8_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10528 = {{4'd0}, _ans_8_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_65 = _GEN_10528 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_67 = {_ans_8_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_69 = _ans_8_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_70 = _ans_8_leadingZeros_T_65 | _ans_8_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10529 = {{2'd0}, _ans_8_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_75 = _GEN_10529 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_77 = {_ans_8_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_79 = _ans_8_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_80 = _ans_8_leadingZeros_T_75 | _ans_8_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10530 = {{1'd0}, _ans_8_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_85 = _GEN_10530 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_87 = {_ans_8_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_89 = _ans_8_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_8_leadingZeros_T_90 = _ans_8_leadingZeros_T_85 | _ans_8_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_8_leadingZeros_T_93 = {_ans_8_leadingZeros_T_49,_ans_8_leadingZeros_T_90,ans_8_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_8_leadingZeros_T_143 = _ans_8_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_144 = _ans_8_leadingZeros_T_93[46] ? 6'h2e : _ans_8_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_145 = _ans_8_leadingZeros_T_93[45] ? 6'h2d : _ans_8_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_146 = _ans_8_leadingZeros_T_93[44] ? 6'h2c : _ans_8_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_147 = _ans_8_leadingZeros_T_93[43] ? 6'h2b : _ans_8_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_148 = _ans_8_leadingZeros_T_93[42] ? 6'h2a : _ans_8_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_149 = _ans_8_leadingZeros_T_93[41] ? 6'h29 : _ans_8_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_150 = _ans_8_leadingZeros_T_93[40] ? 6'h28 : _ans_8_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_151 = _ans_8_leadingZeros_T_93[39] ? 6'h27 : _ans_8_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_152 = _ans_8_leadingZeros_T_93[38] ? 6'h26 : _ans_8_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_153 = _ans_8_leadingZeros_T_93[37] ? 6'h25 : _ans_8_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_154 = _ans_8_leadingZeros_T_93[36] ? 6'h24 : _ans_8_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_155 = _ans_8_leadingZeros_T_93[35] ? 6'h23 : _ans_8_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_156 = _ans_8_leadingZeros_T_93[34] ? 6'h22 : _ans_8_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_157 = _ans_8_leadingZeros_T_93[33] ? 6'h21 : _ans_8_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_158 = _ans_8_leadingZeros_T_93[32] ? 6'h20 : _ans_8_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_159 = _ans_8_leadingZeros_T_93[31] ? 6'h1f : _ans_8_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_160 = _ans_8_leadingZeros_T_93[30] ? 6'h1e : _ans_8_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_161 = _ans_8_leadingZeros_T_93[29] ? 6'h1d : _ans_8_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_162 = _ans_8_leadingZeros_T_93[28] ? 6'h1c : _ans_8_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_163 = _ans_8_leadingZeros_T_93[27] ? 6'h1b : _ans_8_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_164 = _ans_8_leadingZeros_T_93[26] ? 6'h1a : _ans_8_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_165 = _ans_8_leadingZeros_T_93[25] ? 6'h19 : _ans_8_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_166 = _ans_8_leadingZeros_T_93[24] ? 6'h18 : _ans_8_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_167 = _ans_8_leadingZeros_T_93[23] ? 6'h17 : _ans_8_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_168 = _ans_8_leadingZeros_T_93[22] ? 6'h16 : _ans_8_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_169 = _ans_8_leadingZeros_T_93[21] ? 6'h15 : _ans_8_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_170 = _ans_8_leadingZeros_T_93[20] ? 6'h14 : _ans_8_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_171 = _ans_8_leadingZeros_T_93[19] ? 6'h13 : _ans_8_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_172 = _ans_8_leadingZeros_T_93[18] ? 6'h12 : _ans_8_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_173 = _ans_8_leadingZeros_T_93[17] ? 6'h11 : _ans_8_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_174 = _ans_8_leadingZeros_T_93[16] ? 6'h10 : _ans_8_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_175 = _ans_8_leadingZeros_T_93[15] ? 6'hf : _ans_8_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_176 = _ans_8_leadingZeros_T_93[14] ? 6'he : _ans_8_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_177 = _ans_8_leadingZeros_T_93[13] ? 6'hd : _ans_8_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_178 = _ans_8_leadingZeros_T_93[12] ? 6'hc : _ans_8_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_179 = _ans_8_leadingZeros_T_93[11] ? 6'hb : _ans_8_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_180 = _ans_8_leadingZeros_T_93[10] ? 6'ha : _ans_8_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_181 = _ans_8_leadingZeros_T_93[9] ? 6'h9 : _ans_8_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_182 = _ans_8_leadingZeros_T_93[8] ? 6'h8 : _ans_8_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_183 = _ans_8_leadingZeros_T_93[7] ? 6'h7 : _ans_8_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_184 = _ans_8_leadingZeros_T_93[6] ? 6'h6 : _ans_8_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_185 = _ans_8_leadingZeros_T_93[5] ? 6'h5 : _ans_8_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_186 = _ans_8_leadingZeros_T_93[4] ? 6'h4 : _ans_8_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_187 = _ans_8_leadingZeros_T_93[3] ? 6'h3 : _ans_8_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_188 = _ans_8_leadingZeros_T_93[2] ? 6'h2 : _ans_8_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_189 = _ans_8_leadingZeros_T_93[1] ? 6'h1 : _ans_8_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_8_leadingZeros = _ans_8_leadingZeros_T_93[0] ? 6'h0 : _ans_8_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_expRaw_T_1 = 6'h1f - ans_8_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_8_expRaw = ans_8_isZero ? 6'h0 : _ans_8_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_8_shiftAmt_T_2 = ans_8_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_8_shiftAmt = ans_8_expRaw > 6'h3 ? _ans_8_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_8_mantissaRaw_T = ans_8_absClipped >> ans_8_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_8_mantissaRaw = _ans_8_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_8_mantissa = ans_8_expRaw >= 6'h3 ? ans_8_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_8_expAdjusted = ans_8_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_8_exp_T_4 = ans_8_expAdjusted > 7'hf ? 4'hf : ans_8_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_8_exp = ans_8_isZero ? 4'h0 : _ans_8_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_8_fp8 = {ans_8_clippedX[31],ans_8_exp,ans_8_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_9 = {24'h0,linear_bias_9}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_9 = tempSum_9 + biasExtended_9; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_9_sign = sum32_9[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_9_absX_T = ~sum32_9; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_9_absX_T_2 = _ans_9_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_9_absX = ans_9_sign ? _ans_9_absX_T_2 : sum32_9; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_9_shiftedX_T_1 = _GEN_10432 - ans_9_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_9_shiftedX_T_3 = ans_9_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_9_shiftedX = ans_9_sign ? _ans_9_shiftedX_T_1 : _ans_9_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_9_scaledX_T_1 = ans_9_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_9_scaledX = _ans_9_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_9_clippedX_T_2 = ans_9_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_9_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_9_clippedX = ans_9_scaledX > 49'h1c0 ? 49'h1c0 : _ans_9_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_9_absClipped_T_1 = ~ans_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_9_absClipped_T_3 = _ans_9_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_9_absClipped = ans_9_clippedX[31] ? _ans_9_absClipped_T_3 : ans_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_9_isZero = ans_9_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10533 = {{16'd0}, ans_9_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_4 = _GEN_10533 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_6 = {ans_9_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_8 = _ans_9_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_9 = _ans_9_leadingZeros_T_4 | _ans_9_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10534 = {{8'd0}, _ans_9_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_14 = _GEN_10534 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_16 = {_ans_9_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_18 = _ans_9_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_19 = _ans_9_leadingZeros_T_14 | _ans_9_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10535 = {{4'd0}, _ans_9_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_24 = _GEN_10535 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_26 = {_ans_9_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_28 = _ans_9_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_29 = _ans_9_leadingZeros_T_24 | _ans_9_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10536 = {{2'd0}, _ans_9_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_34 = _GEN_10536 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_36 = {_ans_9_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_38 = _ans_9_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_39 = _ans_9_leadingZeros_T_34 | _ans_9_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10537 = {{1'd0}, _ans_9_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_44 = _GEN_10537 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_46 = {_ans_9_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_48 = _ans_9_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_9_leadingZeros_T_49 = _ans_9_leadingZeros_T_44 | _ans_9_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10538 = {{8'd0}, ans_9_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_55 = _GEN_10538 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_57 = {ans_9_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_59 = _ans_9_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_60 = _ans_9_leadingZeros_T_55 | _ans_9_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10539 = {{4'd0}, _ans_9_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_65 = _GEN_10539 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_67 = {_ans_9_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_69 = _ans_9_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_70 = _ans_9_leadingZeros_T_65 | _ans_9_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10540 = {{2'd0}, _ans_9_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_75 = _GEN_10540 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_77 = {_ans_9_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_79 = _ans_9_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_80 = _ans_9_leadingZeros_T_75 | _ans_9_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10541 = {{1'd0}, _ans_9_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_85 = _GEN_10541 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_87 = {_ans_9_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_89 = _ans_9_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_9_leadingZeros_T_90 = _ans_9_leadingZeros_T_85 | _ans_9_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_9_leadingZeros_T_93 = {_ans_9_leadingZeros_T_49,_ans_9_leadingZeros_T_90,ans_9_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_9_leadingZeros_T_143 = _ans_9_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_144 = _ans_9_leadingZeros_T_93[46] ? 6'h2e : _ans_9_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_145 = _ans_9_leadingZeros_T_93[45] ? 6'h2d : _ans_9_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_146 = _ans_9_leadingZeros_T_93[44] ? 6'h2c : _ans_9_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_147 = _ans_9_leadingZeros_T_93[43] ? 6'h2b : _ans_9_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_148 = _ans_9_leadingZeros_T_93[42] ? 6'h2a : _ans_9_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_149 = _ans_9_leadingZeros_T_93[41] ? 6'h29 : _ans_9_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_150 = _ans_9_leadingZeros_T_93[40] ? 6'h28 : _ans_9_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_151 = _ans_9_leadingZeros_T_93[39] ? 6'h27 : _ans_9_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_152 = _ans_9_leadingZeros_T_93[38] ? 6'h26 : _ans_9_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_153 = _ans_9_leadingZeros_T_93[37] ? 6'h25 : _ans_9_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_154 = _ans_9_leadingZeros_T_93[36] ? 6'h24 : _ans_9_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_155 = _ans_9_leadingZeros_T_93[35] ? 6'h23 : _ans_9_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_156 = _ans_9_leadingZeros_T_93[34] ? 6'h22 : _ans_9_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_157 = _ans_9_leadingZeros_T_93[33] ? 6'h21 : _ans_9_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_158 = _ans_9_leadingZeros_T_93[32] ? 6'h20 : _ans_9_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_159 = _ans_9_leadingZeros_T_93[31] ? 6'h1f : _ans_9_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_160 = _ans_9_leadingZeros_T_93[30] ? 6'h1e : _ans_9_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_161 = _ans_9_leadingZeros_T_93[29] ? 6'h1d : _ans_9_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_162 = _ans_9_leadingZeros_T_93[28] ? 6'h1c : _ans_9_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_163 = _ans_9_leadingZeros_T_93[27] ? 6'h1b : _ans_9_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_164 = _ans_9_leadingZeros_T_93[26] ? 6'h1a : _ans_9_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_165 = _ans_9_leadingZeros_T_93[25] ? 6'h19 : _ans_9_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_166 = _ans_9_leadingZeros_T_93[24] ? 6'h18 : _ans_9_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_167 = _ans_9_leadingZeros_T_93[23] ? 6'h17 : _ans_9_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_168 = _ans_9_leadingZeros_T_93[22] ? 6'h16 : _ans_9_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_169 = _ans_9_leadingZeros_T_93[21] ? 6'h15 : _ans_9_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_170 = _ans_9_leadingZeros_T_93[20] ? 6'h14 : _ans_9_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_171 = _ans_9_leadingZeros_T_93[19] ? 6'h13 : _ans_9_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_172 = _ans_9_leadingZeros_T_93[18] ? 6'h12 : _ans_9_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_173 = _ans_9_leadingZeros_T_93[17] ? 6'h11 : _ans_9_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_174 = _ans_9_leadingZeros_T_93[16] ? 6'h10 : _ans_9_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_175 = _ans_9_leadingZeros_T_93[15] ? 6'hf : _ans_9_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_176 = _ans_9_leadingZeros_T_93[14] ? 6'he : _ans_9_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_177 = _ans_9_leadingZeros_T_93[13] ? 6'hd : _ans_9_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_178 = _ans_9_leadingZeros_T_93[12] ? 6'hc : _ans_9_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_179 = _ans_9_leadingZeros_T_93[11] ? 6'hb : _ans_9_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_180 = _ans_9_leadingZeros_T_93[10] ? 6'ha : _ans_9_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_181 = _ans_9_leadingZeros_T_93[9] ? 6'h9 : _ans_9_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_182 = _ans_9_leadingZeros_T_93[8] ? 6'h8 : _ans_9_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_183 = _ans_9_leadingZeros_T_93[7] ? 6'h7 : _ans_9_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_184 = _ans_9_leadingZeros_T_93[6] ? 6'h6 : _ans_9_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_185 = _ans_9_leadingZeros_T_93[5] ? 6'h5 : _ans_9_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_186 = _ans_9_leadingZeros_T_93[4] ? 6'h4 : _ans_9_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_187 = _ans_9_leadingZeros_T_93[3] ? 6'h3 : _ans_9_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_188 = _ans_9_leadingZeros_T_93[2] ? 6'h2 : _ans_9_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_189 = _ans_9_leadingZeros_T_93[1] ? 6'h1 : _ans_9_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_9_leadingZeros = _ans_9_leadingZeros_T_93[0] ? 6'h0 : _ans_9_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_expRaw_T_1 = 6'h1f - ans_9_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_9_expRaw = ans_9_isZero ? 6'h0 : _ans_9_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_9_shiftAmt_T_2 = ans_9_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_9_shiftAmt = ans_9_expRaw > 6'h3 ? _ans_9_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_9_mantissaRaw_T = ans_9_absClipped >> ans_9_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_9_mantissaRaw = _ans_9_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_9_mantissa = ans_9_expRaw >= 6'h3 ? ans_9_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_9_expAdjusted = ans_9_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_9_exp_T_4 = ans_9_expAdjusted > 7'hf ? 4'hf : ans_9_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_9_exp = ans_9_isZero ? 4'h0 : _ans_9_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_9_fp8 = {ans_9_clippedX[31],ans_9_exp,ans_9_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_10 = {24'h0,linear_bias_10}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_10 = tempSum_10 + biasExtended_10; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_10_sign = sum32_10[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_10_absX_T = ~sum32_10; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_10_absX_T_2 = _ans_10_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_10_absX = ans_10_sign ? _ans_10_absX_T_2 : sum32_10; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_10_shiftedX_T_1 = _GEN_10432 - ans_10_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_10_shiftedX_T_3 = ans_10_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_10_shiftedX = ans_10_sign ? _ans_10_shiftedX_T_1 : _ans_10_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_10_scaledX_T_1 = ans_10_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_10_scaledX = _ans_10_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_10_clippedX_T_2 = ans_10_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_10_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_10_clippedX = ans_10_scaledX > 49'h1c0 ? 49'h1c0 : _ans_10_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_10_absClipped_T_1 = ~ans_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_10_absClipped_T_3 = _ans_10_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_10_absClipped = ans_10_clippedX[31] ? _ans_10_absClipped_T_3 : ans_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_10_isZero = ans_10_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10544 = {{16'd0}, ans_10_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_4 = _GEN_10544 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_6 = {ans_10_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_8 = _ans_10_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_9 = _ans_10_leadingZeros_T_4 | _ans_10_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10545 = {{8'd0}, _ans_10_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_14 = _GEN_10545 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_16 = {_ans_10_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_18 = _ans_10_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_19 = _ans_10_leadingZeros_T_14 | _ans_10_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10546 = {{4'd0}, _ans_10_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_24 = _GEN_10546 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_26 = {_ans_10_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_28 = _ans_10_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_29 = _ans_10_leadingZeros_T_24 | _ans_10_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10547 = {{2'd0}, _ans_10_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_34 = _GEN_10547 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_36 = {_ans_10_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_38 = _ans_10_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_39 = _ans_10_leadingZeros_T_34 | _ans_10_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10548 = {{1'd0}, _ans_10_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_44 = _GEN_10548 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_46 = {_ans_10_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_48 = _ans_10_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_10_leadingZeros_T_49 = _ans_10_leadingZeros_T_44 | _ans_10_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10549 = {{8'd0}, ans_10_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_55 = _GEN_10549 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_57 = {ans_10_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_59 = _ans_10_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_60 = _ans_10_leadingZeros_T_55 | _ans_10_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10550 = {{4'd0}, _ans_10_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_65 = _GEN_10550 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_67 = {_ans_10_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_69 = _ans_10_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_70 = _ans_10_leadingZeros_T_65 | _ans_10_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10551 = {{2'd0}, _ans_10_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_75 = _GEN_10551 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_77 = {_ans_10_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_79 = _ans_10_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_80 = _ans_10_leadingZeros_T_75 | _ans_10_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10552 = {{1'd0}, _ans_10_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_85 = _GEN_10552 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_87 = {_ans_10_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_89 = _ans_10_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_10_leadingZeros_T_90 = _ans_10_leadingZeros_T_85 | _ans_10_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_10_leadingZeros_T_93 = {_ans_10_leadingZeros_T_49,_ans_10_leadingZeros_T_90,ans_10_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_10_leadingZeros_T_143 = _ans_10_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_144 = _ans_10_leadingZeros_T_93[46] ? 6'h2e : _ans_10_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_145 = _ans_10_leadingZeros_T_93[45] ? 6'h2d : _ans_10_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_146 = _ans_10_leadingZeros_T_93[44] ? 6'h2c : _ans_10_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_147 = _ans_10_leadingZeros_T_93[43] ? 6'h2b : _ans_10_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_148 = _ans_10_leadingZeros_T_93[42] ? 6'h2a : _ans_10_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_149 = _ans_10_leadingZeros_T_93[41] ? 6'h29 : _ans_10_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_150 = _ans_10_leadingZeros_T_93[40] ? 6'h28 : _ans_10_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_151 = _ans_10_leadingZeros_T_93[39] ? 6'h27 : _ans_10_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_152 = _ans_10_leadingZeros_T_93[38] ? 6'h26 : _ans_10_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_153 = _ans_10_leadingZeros_T_93[37] ? 6'h25 : _ans_10_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_154 = _ans_10_leadingZeros_T_93[36] ? 6'h24 : _ans_10_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_155 = _ans_10_leadingZeros_T_93[35] ? 6'h23 : _ans_10_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_156 = _ans_10_leadingZeros_T_93[34] ? 6'h22 : _ans_10_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_157 = _ans_10_leadingZeros_T_93[33] ? 6'h21 : _ans_10_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_158 = _ans_10_leadingZeros_T_93[32] ? 6'h20 : _ans_10_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_159 = _ans_10_leadingZeros_T_93[31] ? 6'h1f : _ans_10_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_160 = _ans_10_leadingZeros_T_93[30] ? 6'h1e : _ans_10_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_161 = _ans_10_leadingZeros_T_93[29] ? 6'h1d : _ans_10_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_162 = _ans_10_leadingZeros_T_93[28] ? 6'h1c : _ans_10_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_163 = _ans_10_leadingZeros_T_93[27] ? 6'h1b : _ans_10_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_164 = _ans_10_leadingZeros_T_93[26] ? 6'h1a : _ans_10_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_165 = _ans_10_leadingZeros_T_93[25] ? 6'h19 : _ans_10_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_166 = _ans_10_leadingZeros_T_93[24] ? 6'h18 : _ans_10_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_167 = _ans_10_leadingZeros_T_93[23] ? 6'h17 : _ans_10_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_168 = _ans_10_leadingZeros_T_93[22] ? 6'h16 : _ans_10_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_169 = _ans_10_leadingZeros_T_93[21] ? 6'h15 : _ans_10_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_170 = _ans_10_leadingZeros_T_93[20] ? 6'h14 : _ans_10_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_171 = _ans_10_leadingZeros_T_93[19] ? 6'h13 : _ans_10_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_172 = _ans_10_leadingZeros_T_93[18] ? 6'h12 : _ans_10_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_173 = _ans_10_leadingZeros_T_93[17] ? 6'h11 : _ans_10_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_174 = _ans_10_leadingZeros_T_93[16] ? 6'h10 : _ans_10_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_175 = _ans_10_leadingZeros_T_93[15] ? 6'hf : _ans_10_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_176 = _ans_10_leadingZeros_T_93[14] ? 6'he : _ans_10_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_177 = _ans_10_leadingZeros_T_93[13] ? 6'hd : _ans_10_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_178 = _ans_10_leadingZeros_T_93[12] ? 6'hc : _ans_10_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_179 = _ans_10_leadingZeros_T_93[11] ? 6'hb : _ans_10_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_180 = _ans_10_leadingZeros_T_93[10] ? 6'ha : _ans_10_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_181 = _ans_10_leadingZeros_T_93[9] ? 6'h9 : _ans_10_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_182 = _ans_10_leadingZeros_T_93[8] ? 6'h8 : _ans_10_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_183 = _ans_10_leadingZeros_T_93[7] ? 6'h7 : _ans_10_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_184 = _ans_10_leadingZeros_T_93[6] ? 6'h6 : _ans_10_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_185 = _ans_10_leadingZeros_T_93[5] ? 6'h5 : _ans_10_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_186 = _ans_10_leadingZeros_T_93[4] ? 6'h4 : _ans_10_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_187 = _ans_10_leadingZeros_T_93[3] ? 6'h3 : _ans_10_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_188 = _ans_10_leadingZeros_T_93[2] ? 6'h2 : _ans_10_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_189 = _ans_10_leadingZeros_T_93[1] ? 6'h1 : _ans_10_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_10_leadingZeros = _ans_10_leadingZeros_T_93[0] ? 6'h0 : _ans_10_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_expRaw_T_1 = 6'h1f - ans_10_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_10_expRaw = ans_10_isZero ? 6'h0 : _ans_10_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_10_shiftAmt_T_2 = ans_10_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_10_shiftAmt = ans_10_expRaw > 6'h3 ? _ans_10_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_10_mantissaRaw_T = ans_10_absClipped >> ans_10_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_10_mantissaRaw = _ans_10_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_10_mantissa = ans_10_expRaw >= 6'h3 ? ans_10_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_10_expAdjusted = ans_10_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_10_exp_T_4 = ans_10_expAdjusted > 7'hf ? 4'hf : ans_10_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_10_exp = ans_10_isZero ? 4'h0 : _ans_10_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_10_fp8 = {ans_10_clippedX[31],ans_10_exp,ans_10_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_11 = {24'h0,linear_bias_11}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_11 = tempSum_11 + biasExtended_11; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_11_sign = sum32_11[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_11_absX_T = ~sum32_11; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_11_absX_T_2 = _ans_11_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_11_absX = ans_11_sign ? _ans_11_absX_T_2 : sum32_11; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_11_shiftedX_T_1 = _GEN_10432 - ans_11_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_11_shiftedX_T_3 = ans_11_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_11_shiftedX = ans_11_sign ? _ans_11_shiftedX_T_1 : _ans_11_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_11_scaledX_T_1 = ans_11_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_11_scaledX = _ans_11_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_11_clippedX_T_2 = ans_11_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_11_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_11_clippedX = ans_11_scaledX > 49'h1c0 ? 49'h1c0 : _ans_11_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_11_absClipped_T_1 = ~ans_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_11_absClipped_T_3 = _ans_11_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_11_absClipped = ans_11_clippedX[31] ? _ans_11_absClipped_T_3 : ans_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_11_isZero = ans_11_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10555 = {{16'd0}, ans_11_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_4 = _GEN_10555 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_6 = {ans_11_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_8 = _ans_11_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_9 = _ans_11_leadingZeros_T_4 | _ans_11_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10556 = {{8'd0}, _ans_11_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_14 = _GEN_10556 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_16 = {_ans_11_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_18 = _ans_11_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_19 = _ans_11_leadingZeros_T_14 | _ans_11_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10557 = {{4'd0}, _ans_11_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_24 = _GEN_10557 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_26 = {_ans_11_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_28 = _ans_11_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_29 = _ans_11_leadingZeros_T_24 | _ans_11_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10558 = {{2'd0}, _ans_11_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_34 = _GEN_10558 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_36 = {_ans_11_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_38 = _ans_11_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_39 = _ans_11_leadingZeros_T_34 | _ans_11_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10559 = {{1'd0}, _ans_11_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_44 = _GEN_10559 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_46 = {_ans_11_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_48 = _ans_11_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_11_leadingZeros_T_49 = _ans_11_leadingZeros_T_44 | _ans_11_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10560 = {{8'd0}, ans_11_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_55 = _GEN_10560 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_57 = {ans_11_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_59 = _ans_11_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_60 = _ans_11_leadingZeros_T_55 | _ans_11_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10561 = {{4'd0}, _ans_11_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_65 = _GEN_10561 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_67 = {_ans_11_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_69 = _ans_11_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_70 = _ans_11_leadingZeros_T_65 | _ans_11_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10562 = {{2'd0}, _ans_11_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_75 = _GEN_10562 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_77 = {_ans_11_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_79 = _ans_11_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_80 = _ans_11_leadingZeros_T_75 | _ans_11_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10563 = {{1'd0}, _ans_11_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_85 = _GEN_10563 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_87 = {_ans_11_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_89 = _ans_11_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_11_leadingZeros_T_90 = _ans_11_leadingZeros_T_85 | _ans_11_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_11_leadingZeros_T_93 = {_ans_11_leadingZeros_T_49,_ans_11_leadingZeros_T_90,ans_11_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_11_leadingZeros_T_143 = _ans_11_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_144 = _ans_11_leadingZeros_T_93[46] ? 6'h2e : _ans_11_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_145 = _ans_11_leadingZeros_T_93[45] ? 6'h2d : _ans_11_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_146 = _ans_11_leadingZeros_T_93[44] ? 6'h2c : _ans_11_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_147 = _ans_11_leadingZeros_T_93[43] ? 6'h2b : _ans_11_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_148 = _ans_11_leadingZeros_T_93[42] ? 6'h2a : _ans_11_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_149 = _ans_11_leadingZeros_T_93[41] ? 6'h29 : _ans_11_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_150 = _ans_11_leadingZeros_T_93[40] ? 6'h28 : _ans_11_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_151 = _ans_11_leadingZeros_T_93[39] ? 6'h27 : _ans_11_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_152 = _ans_11_leadingZeros_T_93[38] ? 6'h26 : _ans_11_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_153 = _ans_11_leadingZeros_T_93[37] ? 6'h25 : _ans_11_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_154 = _ans_11_leadingZeros_T_93[36] ? 6'h24 : _ans_11_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_155 = _ans_11_leadingZeros_T_93[35] ? 6'h23 : _ans_11_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_156 = _ans_11_leadingZeros_T_93[34] ? 6'h22 : _ans_11_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_157 = _ans_11_leadingZeros_T_93[33] ? 6'h21 : _ans_11_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_158 = _ans_11_leadingZeros_T_93[32] ? 6'h20 : _ans_11_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_159 = _ans_11_leadingZeros_T_93[31] ? 6'h1f : _ans_11_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_160 = _ans_11_leadingZeros_T_93[30] ? 6'h1e : _ans_11_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_161 = _ans_11_leadingZeros_T_93[29] ? 6'h1d : _ans_11_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_162 = _ans_11_leadingZeros_T_93[28] ? 6'h1c : _ans_11_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_163 = _ans_11_leadingZeros_T_93[27] ? 6'h1b : _ans_11_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_164 = _ans_11_leadingZeros_T_93[26] ? 6'h1a : _ans_11_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_165 = _ans_11_leadingZeros_T_93[25] ? 6'h19 : _ans_11_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_166 = _ans_11_leadingZeros_T_93[24] ? 6'h18 : _ans_11_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_167 = _ans_11_leadingZeros_T_93[23] ? 6'h17 : _ans_11_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_168 = _ans_11_leadingZeros_T_93[22] ? 6'h16 : _ans_11_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_169 = _ans_11_leadingZeros_T_93[21] ? 6'h15 : _ans_11_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_170 = _ans_11_leadingZeros_T_93[20] ? 6'h14 : _ans_11_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_171 = _ans_11_leadingZeros_T_93[19] ? 6'h13 : _ans_11_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_172 = _ans_11_leadingZeros_T_93[18] ? 6'h12 : _ans_11_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_173 = _ans_11_leadingZeros_T_93[17] ? 6'h11 : _ans_11_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_174 = _ans_11_leadingZeros_T_93[16] ? 6'h10 : _ans_11_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_175 = _ans_11_leadingZeros_T_93[15] ? 6'hf : _ans_11_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_176 = _ans_11_leadingZeros_T_93[14] ? 6'he : _ans_11_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_177 = _ans_11_leadingZeros_T_93[13] ? 6'hd : _ans_11_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_178 = _ans_11_leadingZeros_T_93[12] ? 6'hc : _ans_11_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_179 = _ans_11_leadingZeros_T_93[11] ? 6'hb : _ans_11_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_180 = _ans_11_leadingZeros_T_93[10] ? 6'ha : _ans_11_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_181 = _ans_11_leadingZeros_T_93[9] ? 6'h9 : _ans_11_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_182 = _ans_11_leadingZeros_T_93[8] ? 6'h8 : _ans_11_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_183 = _ans_11_leadingZeros_T_93[7] ? 6'h7 : _ans_11_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_184 = _ans_11_leadingZeros_T_93[6] ? 6'h6 : _ans_11_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_185 = _ans_11_leadingZeros_T_93[5] ? 6'h5 : _ans_11_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_186 = _ans_11_leadingZeros_T_93[4] ? 6'h4 : _ans_11_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_187 = _ans_11_leadingZeros_T_93[3] ? 6'h3 : _ans_11_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_188 = _ans_11_leadingZeros_T_93[2] ? 6'h2 : _ans_11_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_189 = _ans_11_leadingZeros_T_93[1] ? 6'h1 : _ans_11_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_11_leadingZeros = _ans_11_leadingZeros_T_93[0] ? 6'h0 : _ans_11_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_expRaw_T_1 = 6'h1f - ans_11_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_11_expRaw = ans_11_isZero ? 6'h0 : _ans_11_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_11_shiftAmt_T_2 = ans_11_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_11_shiftAmt = ans_11_expRaw > 6'h3 ? _ans_11_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_11_mantissaRaw_T = ans_11_absClipped >> ans_11_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_11_mantissaRaw = _ans_11_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_11_mantissa = ans_11_expRaw >= 6'h3 ? ans_11_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_11_expAdjusted = ans_11_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_11_exp_T_4 = ans_11_expAdjusted > 7'hf ? 4'hf : ans_11_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_11_exp = ans_11_isZero ? 4'h0 : _ans_11_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_11_fp8 = {ans_11_clippedX[31],ans_11_exp,ans_11_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_12 = {24'h0,linear_bias_12}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_12 = tempSum_12 + biasExtended_12; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_12_sign = sum32_12[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_12_absX_T = ~sum32_12; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_12_absX_T_2 = _ans_12_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_12_absX = ans_12_sign ? _ans_12_absX_T_2 : sum32_12; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_12_shiftedX_T_1 = _GEN_10432 - ans_12_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_12_shiftedX_T_3 = ans_12_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_12_shiftedX = ans_12_sign ? _ans_12_shiftedX_T_1 : _ans_12_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_12_scaledX_T_1 = ans_12_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_12_scaledX = _ans_12_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_12_clippedX_T_2 = ans_12_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_12_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_12_clippedX = ans_12_scaledX > 49'h1c0 ? 49'h1c0 : _ans_12_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_12_absClipped_T_1 = ~ans_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_12_absClipped_T_3 = _ans_12_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_12_absClipped = ans_12_clippedX[31] ? _ans_12_absClipped_T_3 : ans_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_12_isZero = ans_12_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10566 = {{16'd0}, ans_12_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_4 = _GEN_10566 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_6 = {ans_12_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_8 = _ans_12_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_9 = _ans_12_leadingZeros_T_4 | _ans_12_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10567 = {{8'd0}, _ans_12_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_14 = _GEN_10567 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_16 = {_ans_12_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_18 = _ans_12_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_19 = _ans_12_leadingZeros_T_14 | _ans_12_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10568 = {{4'd0}, _ans_12_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_24 = _GEN_10568 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_26 = {_ans_12_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_28 = _ans_12_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_29 = _ans_12_leadingZeros_T_24 | _ans_12_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10569 = {{2'd0}, _ans_12_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_34 = _GEN_10569 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_36 = {_ans_12_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_38 = _ans_12_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_39 = _ans_12_leadingZeros_T_34 | _ans_12_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10570 = {{1'd0}, _ans_12_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_44 = _GEN_10570 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_46 = {_ans_12_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_48 = _ans_12_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_12_leadingZeros_T_49 = _ans_12_leadingZeros_T_44 | _ans_12_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10571 = {{8'd0}, ans_12_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_55 = _GEN_10571 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_57 = {ans_12_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_59 = _ans_12_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_60 = _ans_12_leadingZeros_T_55 | _ans_12_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10572 = {{4'd0}, _ans_12_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_65 = _GEN_10572 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_67 = {_ans_12_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_69 = _ans_12_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_70 = _ans_12_leadingZeros_T_65 | _ans_12_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10573 = {{2'd0}, _ans_12_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_75 = _GEN_10573 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_77 = {_ans_12_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_79 = _ans_12_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_80 = _ans_12_leadingZeros_T_75 | _ans_12_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10574 = {{1'd0}, _ans_12_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_85 = _GEN_10574 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_87 = {_ans_12_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_89 = _ans_12_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_12_leadingZeros_T_90 = _ans_12_leadingZeros_T_85 | _ans_12_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_12_leadingZeros_T_93 = {_ans_12_leadingZeros_T_49,_ans_12_leadingZeros_T_90,ans_12_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_12_leadingZeros_T_143 = _ans_12_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_144 = _ans_12_leadingZeros_T_93[46] ? 6'h2e : _ans_12_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_145 = _ans_12_leadingZeros_T_93[45] ? 6'h2d : _ans_12_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_146 = _ans_12_leadingZeros_T_93[44] ? 6'h2c : _ans_12_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_147 = _ans_12_leadingZeros_T_93[43] ? 6'h2b : _ans_12_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_148 = _ans_12_leadingZeros_T_93[42] ? 6'h2a : _ans_12_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_149 = _ans_12_leadingZeros_T_93[41] ? 6'h29 : _ans_12_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_150 = _ans_12_leadingZeros_T_93[40] ? 6'h28 : _ans_12_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_151 = _ans_12_leadingZeros_T_93[39] ? 6'h27 : _ans_12_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_152 = _ans_12_leadingZeros_T_93[38] ? 6'h26 : _ans_12_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_153 = _ans_12_leadingZeros_T_93[37] ? 6'h25 : _ans_12_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_154 = _ans_12_leadingZeros_T_93[36] ? 6'h24 : _ans_12_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_155 = _ans_12_leadingZeros_T_93[35] ? 6'h23 : _ans_12_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_156 = _ans_12_leadingZeros_T_93[34] ? 6'h22 : _ans_12_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_157 = _ans_12_leadingZeros_T_93[33] ? 6'h21 : _ans_12_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_158 = _ans_12_leadingZeros_T_93[32] ? 6'h20 : _ans_12_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_159 = _ans_12_leadingZeros_T_93[31] ? 6'h1f : _ans_12_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_160 = _ans_12_leadingZeros_T_93[30] ? 6'h1e : _ans_12_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_161 = _ans_12_leadingZeros_T_93[29] ? 6'h1d : _ans_12_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_162 = _ans_12_leadingZeros_T_93[28] ? 6'h1c : _ans_12_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_163 = _ans_12_leadingZeros_T_93[27] ? 6'h1b : _ans_12_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_164 = _ans_12_leadingZeros_T_93[26] ? 6'h1a : _ans_12_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_165 = _ans_12_leadingZeros_T_93[25] ? 6'h19 : _ans_12_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_166 = _ans_12_leadingZeros_T_93[24] ? 6'h18 : _ans_12_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_167 = _ans_12_leadingZeros_T_93[23] ? 6'h17 : _ans_12_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_168 = _ans_12_leadingZeros_T_93[22] ? 6'h16 : _ans_12_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_169 = _ans_12_leadingZeros_T_93[21] ? 6'h15 : _ans_12_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_170 = _ans_12_leadingZeros_T_93[20] ? 6'h14 : _ans_12_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_171 = _ans_12_leadingZeros_T_93[19] ? 6'h13 : _ans_12_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_172 = _ans_12_leadingZeros_T_93[18] ? 6'h12 : _ans_12_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_173 = _ans_12_leadingZeros_T_93[17] ? 6'h11 : _ans_12_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_174 = _ans_12_leadingZeros_T_93[16] ? 6'h10 : _ans_12_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_175 = _ans_12_leadingZeros_T_93[15] ? 6'hf : _ans_12_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_176 = _ans_12_leadingZeros_T_93[14] ? 6'he : _ans_12_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_177 = _ans_12_leadingZeros_T_93[13] ? 6'hd : _ans_12_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_178 = _ans_12_leadingZeros_T_93[12] ? 6'hc : _ans_12_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_179 = _ans_12_leadingZeros_T_93[11] ? 6'hb : _ans_12_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_180 = _ans_12_leadingZeros_T_93[10] ? 6'ha : _ans_12_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_181 = _ans_12_leadingZeros_T_93[9] ? 6'h9 : _ans_12_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_182 = _ans_12_leadingZeros_T_93[8] ? 6'h8 : _ans_12_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_183 = _ans_12_leadingZeros_T_93[7] ? 6'h7 : _ans_12_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_184 = _ans_12_leadingZeros_T_93[6] ? 6'h6 : _ans_12_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_185 = _ans_12_leadingZeros_T_93[5] ? 6'h5 : _ans_12_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_186 = _ans_12_leadingZeros_T_93[4] ? 6'h4 : _ans_12_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_187 = _ans_12_leadingZeros_T_93[3] ? 6'h3 : _ans_12_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_188 = _ans_12_leadingZeros_T_93[2] ? 6'h2 : _ans_12_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_189 = _ans_12_leadingZeros_T_93[1] ? 6'h1 : _ans_12_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_12_leadingZeros = _ans_12_leadingZeros_T_93[0] ? 6'h0 : _ans_12_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_expRaw_T_1 = 6'h1f - ans_12_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_12_expRaw = ans_12_isZero ? 6'h0 : _ans_12_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_12_shiftAmt_T_2 = ans_12_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_12_shiftAmt = ans_12_expRaw > 6'h3 ? _ans_12_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_12_mantissaRaw_T = ans_12_absClipped >> ans_12_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_12_mantissaRaw = _ans_12_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_12_mantissa = ans_12_expRaw >= 6'h3 ? ans_12_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_12_expAdjusted = ans_12_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_12_exp_T_4 = ans_12_expAdjusted > 7'hf ? 4'hf : ans_12_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_12_exp = ans_12_isZero ? 4'h0 : _ans_12_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_12_fp8 = {ans_12_clippedX[31],ans_12_exp,ans_12_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_13 = {24'h0,linear_bias_13}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_13 = tempSum_13 + biasExtended_13; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_13_sign = sum32_13[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_13_absX_T = ~sum32_13; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_13_absX_T_2 = _ans_13_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_13_absX = ans_13_sign ? _ans_13_absX_T_2 : sum32_13; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_13_shiftedX_T_1 = _GEN_10432 - ans_13_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_13_shiftedX_T_3 = ans_13_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_13_shiftedX = ans_13_sign ? _ans_13_shiftedX_T_1 : _ans_13_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_13_scaledX_T_1 = ans_13_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_13_scaledX = _ans_13_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_13_clippedX_T_2 = ans_13_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_13_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_13_clippedX = ans_13_scaledX > 49'h1c0 ? 49'h1c0 : _ans_13_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_13_absClipped_T_1 = ~ans_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_13_absClipped_T_3 = _ans_13_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_13_absClipped = ans_13_clippedX[31] ? _ans_13_absClipped_T_3 : ans_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_13_isZero = ans_13_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10577 = {{16'd0}, ans_13_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_4 = _GEN_10577 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_6 = {ans_13_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_8 = _ans_13_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_9 = _ans_13_leadingZeros_T_4 | _ans_13_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10578 = {{8'd0}, _ans_13_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_14 = _GEN_10578 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_16 = {_ans_13_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_18 = _ans_13_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_19 = _ans_13_leadingZeros_T_14 | _ans_13_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10579 = {{4'd0}, _ans_13_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_24 = _GEN_10579 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_26 = {_ans_13_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_28 = _ans_13_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_29 = _ans_13_leadingZeros_T_24 | _ans_13_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10580 = {{2'd0}, _ans_13_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_34 = _GEN_10580 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_36 = {_ans_13_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_38 = _ans_13_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_39 = _ans_13_leadingZeros_T_34 | _ans_13_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10581 = {{1'd0}, _ans_13_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_44 = _GEN_10581 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_46 = {_ans_13_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_48 = _ans_13_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_13_leadingZeros_T_49 = _ans_13_leadingZeros_T_44 | _ans_13_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10582 = {{8'd0}, ans_13_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_55 = _GEN_10582 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_57 = {ans_13_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_59 = _ans_13_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_60 = _ans_13_leadingZeros_T_55 | _ans_13_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10583 = {{4'd0}, _ans_13_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_65 = _GEN_10583 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_67 = {_ans_13_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_69 = _ans_13_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_70 = _ans_13_leadingZeros_T_65 | _ans_13_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10584 = {{2'd0}, _ans_13_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_75 = _GEN_10584 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_77 = {_ans_13_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_79 = _ans_13_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_80 = _ans_13_leadingZeros_T_75 | _ans_13_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10585 = {{1'd0}, _ans_13_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_85 = _GEN_10585 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_87 = {_ans_13_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_89 = _ans_13_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_13_leadingZeros_T_90 = _ans_13_leadingZeros_T_85 | _ans_13_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_13_leadingZeros_T_93 = {_ans_13_leadingZeros_T_49,_ans_13_leadingZeros_T_90,ans_13_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_13_leadingZeros_T_143 = _ans_13_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_144 = _ans_13_leadingZeros_T_93[46] ? 6'h2e : _ans_13_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_145 = _ans_13_leadingZeros_T_93[45] ? 6'h2d : _ans_13_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_146 = _ans_13_leadingZeros_T_93[44] ? 6'h2c : _ans_13_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_147 = _ans_13_leadingZeros_T_93[43] ? 6'h2b : _ans_13_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_148 = _ans_13_leadingZeros_T_93[42] ? 6'h2a : _ans_13_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_149 = _ans_13_leadingZeros_T_93[41] ? 6'h29 : _ans_13_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_150 = _ans_13_leadingZeros_T_93[40] ? 6'h28 : _ans_13_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_151 = _ans_13_leadingZeros_T_93[39] ? 6'h27 : _ans_13_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_152 = _ans_13_leadingZeros_T_93[38] ? 6'h26 : _ans_13_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_153 = _ans_13_leadingZeros_T_93[37] ? 6'h25 : _ans_13_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_154 = _ans_13_leadingZeros_T_93[36] ? 6'h24 : _ans_13_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_155 = _ans_13_leadingZeros_T_93[35] ? 6'h23 : _ans_13_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_156 = _ans_13_leadingZeros_T_93[34] ? 6'h22 : _ans_13_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_157 = _ans_13_leadingZeros_T_93[33] ? 6'h21 : _ans_13_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_158 = _ans_13_leadingZeros_T_93[32] ? 6'h20 : _ans_13_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_159 = _ans_13_leadingZeros_T_93[31] ? 6'h1f : _ans_13_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_160 = _ans_13_leadingZeros_T_93[30] ? 6'h1e : _ans_13_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_161 = _ans_13_leadingZeros_T_93[29] ? 6'h1d : _ans_13_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_162 = _ans_13_leadingZeros_T_93[28] ? 6'h1c : _ans_13_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_163 = _ans_13_leadingZeros_T_93[27] ? 6'h1b : _ans_13_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_164 = _ans_13_leadingZeros_T_93[26] ? 6'h1a : _ans_13_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_165 = _ans_13_leadingZeros_T_93[25] ? 6'h19 : _ans_13_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_166 = _ans_13_leadingZeros_T_93[24] ? 6'h18 : _ans_13_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_167 = _ans_13_leadingZeros_T_93[23] ? 6'h17 : _ans_13_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_168 = _ans_13_leadingZeros_T_93[22] ? 6'h16 : _ans_13_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_169 = _ans_13_leadingZeros_T_93[21] ? 6'h15 : _ans_13_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_170 = _ans_13_leadingZeros_T_93[20] ? 6'h14 : _ans_13_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_171 = _ans_13_leadingZeros_T_93[19] ? 6'h13 : _ans_13_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_172 = _ans_13_leadingZeros_T_93[18] ? 6'h12 : _ans_13_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_173 = _ans_13_leadingZeros_T_93[17] ? 6'h11 : _ans_13_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_174 = _ans_13_leadingZeros_T_93[16] ? 6'h10 : _ans_13_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_175 = _ans_13_leadingZeros_T_93[15] ? 6'hf : _ans_13_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_176 = _ans_13_leadingZeros_T_93[14] ? 6'he : _ans_13_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_177 = _ans_13_leadingZeros_T_93[13] ? 6'hd : _ans_13_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_178 = _ans_13_leadingZeros_T_93[12] ? 6'hc : _ans_13_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_179 = _ans_13_leadingZeros_T_93[11] ? 6'hb : _ans_13_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_180 = _ans_13_leadingZeros_T_93[10] ? 6'ha : _ans_13_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_181 = _ans_13_leadingZeros_T_93[9] ? 6'h9 : _ans_13_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_182 = _ans_13_leadingZeros_T_93[8] ? 6'h8 : _ans_13_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_183 = _ans_13_leadingZeros_T_93[7] ? 6'h7 : _ans_13_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_184 = _ans_13_leadingZeros_T_93[6] ? 6'h6 : _ans_13_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_185 = _ans_13_leadingZeros_T_93[5] ? 6'h5 : _ans_13_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_186 = _ans_13_leadingZeros_T_93[4] ? 6'h4 : _ans_13_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_187 = _ans_13_leadingZeros_T_93[3] ? 6'h3 : _ans_13_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_188 = _ans_13_leadingZeros_T_93[2] ? 6'h2 : _ans_13_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_189 = _ans_13_leadingZeros_T_93[1] ? 6'h1 : _ans_13_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_13_leadingZeros = _ans_13_leadingZeros_T_93[0] ? 6'h0 : _ans_13_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_expRaw_T_1 = 6'h1f - ans_13_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_13_expRaw = ans_13_isZero ? 6'h0 : _ans_13_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_13_shiftAmt_T_2 = ans_13_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_13_shiftAmt = ans_13_expRaw > 6'h3 ? _ans_13_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_13_mantissaRaw_T = ans_13_absClipped >> ans_13_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_13_mantissaRaw = _ans_13_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_13_mantissa = ans_13_expRaw >= 6'h3 ? ans_13_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_13_expAdjusted = ans_13_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_13_exp_T_4 = ans_13_expAdjusted > 7'hf ? 4'hf : ans_13_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_13_exp = ans_13_isZero ? 4'h0 : _ans_13_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_13_fp8 = {ans_13_clippedX[31],ans_13_exp,ans_13_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_14 = {24'h0,linear_bias_14}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_14 = tempSum_14 + biasExtended_14; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_14_sign = sum32_14[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_14_absX_T = ~sum32_14; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_14_absX_T_2 = _ans_14_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_14_absX = ans_14_sign ? _ans_14_absX_T_2 : sum32_14; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_14_shiftedX_T_1 = _GEN_10432 - ans_14_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_14_shiftedX_T_3 = ans_14_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_14_shiftedX = ans_14_sign ? _ans_14_shiftedX_T_1 : _ans_14_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_14_scaledX_T_1 = ans_14_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_14_scaledX = _ans_14_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_14_clippedX_T_2 = ans_14_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_14_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_14_clippedX = ans_14_scaledX > 49'h1c0 ? 49'h1c0 : _ans_14_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_14_absClipped_T_1 = ~ans_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_14_absClipped_T_3 = _ans_14_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_14_absClipped = ans_14_clippedX[31] ? _ans_14_absClipped_T_3 : ans_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_14_isZero = ans_14_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10588 = {{16'd0}, ans_14_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_4 = _GEN_10588 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_6 = {ans_14_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_8 = _ans_14_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_9 = _ans_14_leadingZeros_T_4 | _ans_14_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10589 = {{8'd0}, _ans_14_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_14 = _GEN_10589 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_16 = {_ans_14_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_18 = _ans_14_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_19 = _ans_14_leadingZeros_T_14 | _ans_14_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10590 = {{4'd0}, _ans_14_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_24 = _GEN_10590 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_26 = {_ans_14_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_28 = _ans_14_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_29 = _ans_14_leadingZeros_T_24 | _ans_14_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10591 = {{2'd0}, _ans_14_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_34 = _GEN_10591 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_36 = {_ans_14_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_38 = _ans_14_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_39 = _ans_14_leadingZeros_T_34 | _ans_14_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10592 = {{1'd0}, _ans_14_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_44 = _GEN_10592 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_46 = {_ans_14_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_48 = _ans_14_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_14_leadingZeros_T_49 = _ans_14_leadingZeros_T_44 | _ans_14_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10593 = {{8'd0}, ans_14_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_55 = _GEN_10593 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_57 = {ans_14_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_59 = _ans_14_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_60 = _ans_14_leadingZeros_T_55 | _ans_14_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10594 = {{4'd0}, _ans_14_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_65 = _GEN_10594 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_67 = {_ans_14_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_69 = _ans_14_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_70 = _ans_14_leadingZeros_T_65 | _ans_14_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10595 = {{2'd0}, _ans_14_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_75 = _GEN_10595 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_77 = {_ans_14_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_79 = _ans_14_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_80 = _ans_14_leadingZeros_T_75 | _ans_14_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10596 = {{1'd0}, _ans_14_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_85 = _GEN_10596 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_87 = {_ans_14_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_89 = _ans_14_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_14_leadingZeros_T_90 = _ans_14_leadingZeros_T_85 | _ans_14_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_14_leadingZeros_T_93 = {_ans_14_leadingZeros_T_49,_ans_14_leadingZeros_T_90,ans_14_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_14_leadingZeros_T_143 = _ans_14_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_144 = _ans_14_leadingZeros_T_93[46] ? 6'h2e : _ans_14_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_145 = _ans_14_leadingZeros_T_93[45] ? 6'h2d : _ans_14_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_146 = _ans_14_leadingZeros_T_93[44] ? 6'h2c : _ans_14_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_147 = _ans_14_leadingZeros_T_93[43] ? 6'h2b : _ans_14_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_148 = _ans_14_leadingZeros_T_93[42] ? 6'h2a : _ans_14_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_149 = _ans_14_leadingZeros_T_93[41] ? 6'h29 : _ans_14_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_150 = _ans_14_leadingZeros_T_93[40] ? 6'h28 : _ans_14_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_151 = _ans_14_leadingZeros_T_93[39] ? 6'h27 : _ans_14_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_152 = _ans_14_leadingZeros_T_93[38] ? 6'h26 : _ans_14_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_153 = _ans_14_leadingZeros_T_93[37] ? 6'h25 : _ans_14_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_154 = _ans_14_leadingZeros_T_93[36] ? 6'h24 : _ans_14_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_155 = _ans_14_leadingZeros_T_93[35] ? 6'h23 : _ans_14_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_156 = _ans_14_leadingZeros_T_93[34] ? 6'h22 : _ans_14_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_157 = _ans_14_leadingZeros_T_93[33] ? 6'h21 : _ans_14_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_158 = _ans_14_leadingZeros_T_93[32] ? 6'h20 : _ans_14_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_159 = _ans_14_leadingZeros_T_93[31] ? 6'h1f : _ans_14_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_160 = _ans_14_leadingZeros_T_93[30] ? 6'h1e : _ans_14_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_161 = _ans_14_leadingZeros_T_93[29] ? 6'h1d : _ans_14_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_162 = _ans_14_leadingZeros_T_93[28] ? 6'h1c : _ans_14_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_163 = _ans_14_leadingZeros_T_93[27] ? 6'h1b : _ans_14_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_164 = _ans_14_leadingZeros_T_93[26] ? 6'h1a : _ans_14_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_165 = _ans_14_leadingZeros_T_93[25] ? 6'h19 : _ans_14_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_166 = _ans_14_leadingZeros_T_93[24] ? 6'h18 : _ans_14_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_167 = _ans_14_leadingZeros_T_93[23] ? 6'h17 : _ans_14_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_168 = _ans_14_leadingZeros_T_93[22] ? 6'h16 : _ans_14_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_169 = _ans_14_leadingZeros_T_93[21] ? 6'h15 : _ans_14_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_170 = _ans_14_leadingZeros_T_93[20] ? 6'h14 : _ans_14_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_171 = _ans_14_leadingZeros_T_93[19] ? 6'h13 : _ans_14_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_172 = _ans_14_leadingZeros_T_93[18] ? 6'h12 : _ans_14_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_173 = _ans_14_leadingZeros_T_93[17] ? 6'h11 : _ans_14_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_174 = _ans_14_leadingZeros_T_93[16] ? 6'h10 : _ans_14_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_175 = _ans_14_leadingZeros_T_93[15] ? 6'hf : _ans_14_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_176 = _ans_14_leadingZeros_T_93[14] ? 6'he : _ans_14_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_177 = _ans_14_leadingZeros_T_93[13] ? 6'hd : _ans_14_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_178 = _ans_14_leadingZeros_T_93[12] ? 6'hc : _ans_14_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_179 = _ans_14_leadingZeros_T_93[11] ? 6'hb : _ans_14_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_180 = _ans_14_leadingZeros_T_93[10] ? 6'ha : _ans_14_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_181 = _ans_14_leadingZeros_T_93[9] ? 6'h9 : _ans_14_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_182 = _ans_14_leadingZeros_T_93[8] ? 6'h8 : _ans_14_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_183 = _ans_14_leadingZeros_T_93[7] ? 6'h7 : _ans_14_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_184 = _ans_14_leadingZeros_T_93[6] ? 6'h6 : _ans_14_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_185 = _ans_14_leadingZeros_T_93[5] ? 6'h5 : _ans_14_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_186 = _ans_14_leadingZeros_T_93[4] ? 6'h4 : _ans_14_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_187 = _ans_14_leadingZeros_T_93[3] ? 6'h3 : _ans_14_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_188 = _ans_14_leadingZeros_T_93[2] ? 6'h2 : _ans_14_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_189 = _ans_14_leadingZeros_T_93[1] ? 6'h1 : _ans_14_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_14_leadingZeros = _ans_14_leadingZeros_T_93[0] ? 6'h0 : _ans_14_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_expRaw_T_1 = 6'h1f - ans_14_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_14_expRaw = ans_14_isZero ? 6'h0 : _ans_14_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_14_shiftAmt_T_2 = ans_14_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_14_shiftAmt = ans_14_expRaw > 6'h3 ? _ans_14_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_14_mantissaRaw_T = ans_14_absClipped >> ans_14_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_14_mantissaRaw = _ans_14_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_14_mantissa = ans_14_expRaw >= 6'h3 ? ans_14_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_14_expAdjusted = ans_14_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_14_exp_T_4 = ans_14_expAdjusted > 7'hf ? 4'hf : ans_14_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_14_exp = ans_14_isZero ? 4'h0 : _ans_14_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_14_fp8 = {ans_14_clippedX[31],ans_14_exp,ans_14_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_15 = {24'h0,linear_bias_15}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_15 = tempSum_15 + biasExtended_15; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_15_sign = sum32_15[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_15_absX_T = ~sum32_15; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_15_absX_T_2 = _ans_15_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_15_absX = ans_15_sign ? _ans_15_absX_T_2 : sum32_15; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_15_shiftedX_T_1 = _GEN_10432 - ans_15_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_15_shiftedX_T_3 = ans_15_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_15_shiftedX = ans_15_sign ? _ans_15_shiftedX_T_1 : _ans_15_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_15_scaledX_T_1 = ans_15_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_15_scaledX = _ans_15_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_15_clippedX_T_2 = ans_15_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_15_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_15_clippedX = ans_15_scaledX > 49'h1c0 ? 49'h1c0 : _ans_15_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_15_absClipped_T_1 = ~ans_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_15_absClipped_T_3 = _ans_15_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_15_absClipped = ans_15_clippedX[31] ? _ans_15_absClipped_T_3 : ans_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_15_isZero = ans_15_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10599 = {{16'd0}, ans_15_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_4 = _GEN_10599 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_6 = {ans_15_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_8 = _ans_15_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_9 = _ans_15_leadingZeros_T_4 | _ans_15_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10600 = {{8'd0}, _ans_15_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_14 = _GEN_10600 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_16 = {_ans_15_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_18 = _ans_15_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_19 = _ans_15_leadingZeros_T_14 | _ans_15_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10601 = {{4'd0}, _ans_15_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_24 = _GEN_10601 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_26 = {_ans_15_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_28 = _ans_15_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_29 = _ans_15_leadingZeros_T_24 | _ans_15_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10602 = {{2'd0}, _ans_15_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_34 = _GEN_10602 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_36 = {_ans_15_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_38 = _ans_15_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_39 = _ans_15_leadingZeros_T_34 | _ans_15_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10603 = {{1'd0}, _ans_15_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_44 = _GEN_10603 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_46 = {_ans_15_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_48 = _ans_15_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_15_leadingZeros_T_49 = _ans_15_leadingZeros_T_44 | _ans_15_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10604 = {{8'd0}, ans_15_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_55 = _GEN_10604 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_57 = {ans_15_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_59 = _ans_15_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_60 = _ans_15_leadingZeros_T_55 | _ans_15_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10605 = {{4'd0}, _ans_15_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_65 = _GEN_10605 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_67 = {_ans_15_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_69 = _ans_15_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_70 = _ans_15_leadingZeros_T_65 | _ans_15_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10606 = {{2'd0}, _ans_15_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_75 = _GEN_10606 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_77 = {_ans_15_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_79 = _ans_15_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_80 = _ans_15_leadingZeros_T_75 | _ans_15_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10607 = {{1'd0}, _ans_15_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_85 = _GEN_10607 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_87 = {_ans_15_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_89 = _ans_15_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_15_leadingZeros_T_90 = _ans_15_leadingZeros_T_85 | _ans_15_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_15_leadingZeros_T_93 = {_ans_15_leadingZeros_T_49,_ans_15_leadingZeros_T_90,ans_15_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_15_leadingZeros_T_143 = _ans_15_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_144 = _ans_15_leadingZeros_T_93[46] ? 6'h2e : _ans_15_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_145 = _ans_15_leadingZeros_T_93[45] ? 6'h2d : _ans_15_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_146 = _ans_15_leadingZeros_T_93[44] ? 6'h2c : _ans_15_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_147 = _ans_15_leadingZeros_T_93[43] ? 6'h2b : _ans_15_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_148 = _ans_15_leadingZeros_T_93[42] ? 6'h2a : _ans_15_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_149 = _ans_15_leadingZeros_T_93[41] ? 6'h29 : _ans_15_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_150 = _ans_15_leadingZeros_T_93[40] ? 6'h28 : _ans_15_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_151 = _ans_15_leadingZeros_T_93[39] ? 6'h27 : _ans_15_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_152 = _ans_15_leadingZeros_T_93[38] ? 6'h26 : _ans_15_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_153 = _ans_15_leadingZeros_T_93[37] ? 6'h25 : _ans_15_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_154 = _ans_15_leadingZeros_T_93[36] ? 6'h24 : _ans_15_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_155 = _ans_15_leadingZeros_T_93[35] ? 6'h23 : _ans_15_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_156 = _ans_15_leadingZeros_T_93[34] ? 6'h22 : _ans_15_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_157 = _ans_15_leadingZeros_T_93[33] ? 6'h21 : _ans_15_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_158 = _ans_15_leadingZeros_T_93[32] ? 6'h20 : _ans_15_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_159 = _ans_15_leadingZeros_T_93[31] ? 6'h1f : _ans_15_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_160 = _ans_15_leadingZeros_T_93[30] ? 6'h1e : _ans_15_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_161 = _ans_15_leadingZeros_T_93[29] ? 6'h1d : _ans_15_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_162 = _ans_15_leadingZeros_T_93[28] ? 6'h1c : _ans_15_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_163 = _ans_15_leadingZeros_T_93[27] ? 6'h1b : _ans_15_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_164 = _ans_15_leadingZeros_T_93[26] ? 6'h1a : _ans_15_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_165 = _ans_15_leadingZeros_T_93[25] ? 6'h19 : _ans_15_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_166 = _ans_15_leadingZeros_T_93[24] ? 6'h18 : _ans_15_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_167 = _ans_15_leadingZeros_T_93[23] ? 6'h17 : _ans_15_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_168 = _ans_15_leadingZeros_T_93[22] ? 6'h16 : _ans_15_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_169 = _ans_15_leadingZeros_T_93[21] ? 6'h15 : _ans_15_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_170 = _ans_15_leadingZeros_T_93[20] ? 6'h14 : _ans_15_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_171 = _ans_15_leadingZeros_T_93[19] ? 6'h13 : _ans_15_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_172 = _ans_15_leadingZeros_T_93[18] ? 6'h12 : _ans_15_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_173 = _ans_15_leadingZeros_T_93[17] ? 6'h11 : _ans_15_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_174 = _ans_15_leadingZeros_T_93[16] ? 6'h10 : _ans_15_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_175 = _ans_15_leadingZeros_T_93[15] ? 6'hf : _ans_15_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_176 = _ans_15_leadingZeros_T_93[14] ? 6'he : _ans_15_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_177 = _ans_15_leadingZeros_T_93[13] ? 6'hd : _ans_15_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_178 = _ans_15_leadingZeros_T_93[12] ? 6'hc : _ans_15_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_179 = _ans_15_leadingZeros_T_93[11] ? 6'hb : _ans_15_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_180 = _ans_15_leadingZeros_T_93[10] ? 6'ha : _ans_15_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_181 = _ans_15_leadingZeros_T_93[9] ? 6'h9 : _ans_15_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_182 = _ans_15_leadingZeros_T_93[8] ? 6'h8 : _ans_15_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_183 = _ans_15_leadingZeros_T_93[7] ? 6'h7 : _ans_15_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_184 = _ans_15_leadingZeros_T_93[6] ? 6'h6 : _ans_15_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_185 = _ans_15_leadingZeros_T_93[5] ? 6'h5 : _ans_15_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_186 = _ans_15_leadingZeros_T_93[4] ? 6'h4 : _ans_15_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_187 = _ans_15_leadingZeros_T_93[3] ? 6'h3 : _ans_15_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_188 = _ans_15_leadingZeros_T_93[2] ? 6'h2 : _ans_15_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_189 = _ans_15_leadingZeros_T_93[1] ? 6'h1 : _ans_15_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_15_leadingZeros = _ans_15_leadingZeros_T_93[0] ? 6'h0 : _ans_15_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_expRaw_T_1 = 6'h1f - ans_15_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_15_expRaw = ans_15_isZero ? 6'h0 : _ans_15_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_15_shiftAmt_T_2 = ans_15_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_15_shiftAmt = ans_15_expRaw > 6'h3 ? _ans_15_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_15_mantissaRaw_T = ans_15_absClipped >> ans_15_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_15_mantissaRaw = _ans_15_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_15_mantissa = ans_15_expRaw >= 6'h3 ? ans_15_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_15_expAdjusted = ans_15_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_15_exp_T_4 = ans_15_expAdjusted > 7'hf ? 4'hf : ans_15_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_15_exp = ans_15_isZero ? 4'h0 : _ans_15_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_15_fp8 = {ans_15_clippedX[31],ans_15_exp,ans_15_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_16 = {24'h0,linear_bias_16}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_16 = tempSum_16 + biasExtended_16; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_16_sign = sum32_16[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_16_absX_T = ~sum32_16; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_16_absX_T_2 = _ans_16_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_16_absX = ans_16_sign ? _ans_16_absX_T_2 : sum32_16; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_16_shiftedX_T_1 = _GEN_10432 - ans_16_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_16_shiftedX_T_3 = ans_16_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_16_shiftedX = ans_16_sign ? _ans_16_shiftedX_T_1 : _ans_16_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_16_scaledX_T_1 = ans_16_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_16_scaledX = _ans_16_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_16_clippedX_T_2 = ans_16_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_16_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_16_clippedX = ans_16_scaledX > 49'h1c0 ? 49'h1c0 : _ans_16_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_16_absClipped_T_1 = ~ans_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_16_absClipped_T_3 = _ans_16_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_16_absClipped = ans_16_clippedX[31] ? _ans_16_absClipped_T_3 : ans_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_16_isZero = ans_16_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10610 = {{16'd0}, ans_16_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_4 = _GEN_10610 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_6 = {ans_16_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_8 = _ans_16_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_9 = _ans_16_leadingZeros_T_4 | _ans_16_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10611 = {{8'd0}, _ans_16_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_14 = _GEN_10611 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_16 = {_ans_16_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_18 = _ans_16_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_19 = _ans_16_leadingZeros_T_14 | _ans_16_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10612 = {{4'd0}, _ans_16_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_24 = _GEN_10612 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_26 = {_ans_16_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_28 = _ans_16_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_29 = _ans_16_leadingZeros_T_24 | _ans_16_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10613 = {{2'd0}, _ans_16_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_34 = _GEN_10613 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_36 = {_ans_16_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_38 = _ans_16_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_39 = _ans_16_leadingZeros_T_34 | _ans_16_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10614 = {{1'd0}, _ans_16_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_44 = _GEN_10614 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_46 = {_ans_16_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_48 = _ans_16_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_16_leadingZeros_T_49 = _ans_16_leadingZeros_T_44 | _ans_16_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10615 = {{8'd0}, ans_16_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_55 = _GEN_10615 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_57 = {ans_16_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_59 = _ans_16_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_60 = _ans_16_leadingZeros_T_55 | _ans_16_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10616 = {{4'd0}, _ans_16_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_65 = _GEN_10616 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_67 = {_ans_16_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_69 = _ans_16_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_70 = _ans_16_leadingZeros_T_65 | _ans_16_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10617 = {{2'd0}, _ans_16_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_75 = _GEN_10617 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_77 = {_ans_16_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_79 = _ans_16_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_80 = _ans_16_leadingZeros_T_75 | _ans_16_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10618 = {{1'd0}, _ans_16_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_85 = _GEN_10618 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_87 = {_ans_16_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_89 = _ans_16_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_16_leadingZeros_T_90 = _ans_16_leadingZeros_T_85 | _ans_16_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_16_leadingZeros_T_93 = {_ans_16_leadingZeros_T_49,_ans_16_leadingZeros_T_90,ans_16_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_16_leadingZeros_T_143 = _ans_16_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_144 = _ans_16_leadingZeros_T_93[46] ? 6'h2e : _ans_16_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_145 = _ans_16_leadingZeros_T_93[45] ? 6'h2d : _ans_16_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_146 = _ans_16_leadingZeros_T_93[44] ? 6'h2c : _ans_16_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_147 = _ans_16_leadingZeros_T_93[43] ? 6'h2b : _ans_16_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_148 = _ans_16_leadingZeros_T_93[42] ? 6'h2a : _ans_16_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_149 = _ans_16_leadingZeros_T_93[41] ? 6'h29 : _ans_16_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_150 = _ans_16_leadingZeros_T_93[40] ? 6'h28 : _ans_16_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_151 = _ans_16_leadingZeros_T_93[39] ? 6'h27 : _ans_16_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_152 = _ans_16_leadingZeros_T_93[38] ? 6'h26 : _ans_16_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_153 = _ans_16_leadingZeros_T_93[37] ? 6'h25 : _ans_16_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_154 = _ans_16_leadingZeros_T_93[36] ? 6'h24 : _ans_16_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_155 = _ans_16_leadingZeros_T_93[35] ? 6'h23 : _ans_16_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_156 = _ans_16_leadingZeros_T_93[34] ? 6'h22 : _ans_16_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_157 = _ans_16_leadingZeros_T_93[33] ? 6'h21 : _ans_16_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_158 = _ans_16_leadingZeros_T_93[32] ? 6'h20 : _ans_16_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_159 = _ans_16_leadingZeros_T_93[31] ? 6'h1f : _ans_16_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_160 = _ans_16_leadingZeros_T_93[30] ? 6'h1e : _ans_16_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_161 = _ans_16_leadingZeros_T_93[29] ? 6'h1d : _ans_16_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_162 = _ans_16_leadingZeros_T_93[28] ? 6'h1c : _ans_16_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_163 = _ans_16_leadingZeros_T_93[27] ? 6'h1b : _ans_16_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_164 = _ans_16_leadingZeros_T_93[26] ? 6'h1a : _ans_16_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_165 = _ans_16_leadingZeros_T_93[25] ? 6'h19 : _ans_16_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_166 = _ans_16_leadingZeros_T_93[24] ? 6'h18 : _ans_16_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_167 = _ans_16_leadingZeros_T_93[23] ? 6'h17 : _ans_16_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_168 = _ans_16_leadingZeros_T_93[22] ? 6'h16 : _ans_16_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_169 = _ans_16_leadingZeros_T_93[21] ? 6'h15 : _ans_16_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_170 = _ans_16_leadingZeros_T_93[20] ? 6'h14 : _ans_16_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_171 = _ans_16_leadingZeros_T_93[19] ? 6'h13 : _ans_16_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_172 = _ans_16_leadingZeros_T_93[18] ? 6'h12 : _ans_16_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_173 = _ans_16_leadingZeros_T_93[17] ? 6'h11 : _ans_16_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_174 = _ans_16_leadingZeros_T_93[16] ? 6'h10 : _ans_16_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_175 = _ans_16_leadingZeros_T_93[15] ? 6'hf : _ans_16_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_176 = _ans_16_leadingZeros_T_93[14] ? 6'he : _ans_16_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_177 = _ans_16_leadingZeros_T_93[13] ? 6'hd : _ans_16_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_178 = _ans_16_leadingZeros_T_93[12] ? 6'hc : _ans_16_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_179 = _ans_16_leadingZeros_T_93[11] ? 6'hb : _ans_16_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_180 = _ans_16_leadingZeros_T_93[10] ? 6'ha : _ans_16_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_181 = _ans_16_leadingZeros_T_93[9] ? 6'h9 : _ans_16_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_182 = _ans_16_leadingZeros_T_93[8] ? 6'h8 : _ans_16_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_183 = _ans_16_leadingZeros_T_93[7] ? 6'h7 : _ans_16_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_184 = _ans_16_leadingZeros_T_93[6] ? 6'h6 : _ans_16_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_185 = _ans_16_leadingZeros_T_93[5] ? 6'h5 : _ans_16_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_186 = _ans_16_leadingZeros_T_93[4] ? 6'h4 : _ans_16_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_187 = _ans_16_leadingZeros_T_93[3] ? 6'h3 : _ans_16_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_188 = _ans_16_leadingZeros_T_93[2] ? 6'h2 : _ans_16_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_189 = _ans_16_leadingZeros_T_93[1] ? 6'h1 : _ans_16_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_16_leadingZeros = _ans_16_leadingZeros_T_93[0] ? 6'h0 : _ans_16_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_expRaw_T_1 = 6'h1f - ans_16_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_16_expRaw = ans_16_isZero ? 6'h0 : _ans_16_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_16_shiftAmt_T_2 = ans_16_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_16_shiftAmt = ans_16_expRaw > 6'h3 ? _ans_16_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_16_mantissaRaw_T = ans_16_absClipped >> ans_16_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_16_mantissaRaw = _ans_16_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_16_mantissa = ans_16_expRaw >= 6'h3 ? ans_16_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_16_expAdjusted = ans_16_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_16_exp_T_4 = ans_16_expAdjusted > 7'hf ? 4'hf : ans_16_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_16_exp = ans_16_isZero ? 4'h0 : _ans_16_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_16_fp8 = {ans_16_clippedX[31],ans_16_exp,ans_16_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_17 = {24'h0,linear_bias_17}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_17 = tempSum_17 + biasExtended_17; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_17_sign = sum32_17[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_17_absX_T = ~sum32_17; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_17_absX_T_2 = _ans_17_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_17_absX = ans_17_sign ? _ans_17_absX_T_2 : sum32_17; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_17_shiftedX_T_1 = _GEN_10432 - ans_17_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_17_shiftedX_T_3 = ans_17_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_17_shiftedX = ans_17_sign ? _ans_17_shiftedX_T_1 : _ans_17_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_17_scaledX_T_1 = ans_17_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_17_scaledX = _ans_17_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_17_clippedX_T_2 = ans_17_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_17_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_17_clippedX = ans_17_scaledX > 49'h1c0 ? 49'h1c0 : _ans_17_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_17_absClipped_T_1 = ~ans_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_17_absClipped_T_3 = _ans_17_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_17_absClipped = ans_17_clippedX[31] ? _ans_17_absClipped_T_3 : ans_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_17_isZero = ans_17_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10621 = {{16'd0}, ans_17_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_4 = _GEN_10621 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_6 = {ans_17_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_8 = _ans_17_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_9 = _ans_17_leadingZeros_T_4 | _ans_17_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10622 = {{8'd0}, _ans_17_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_14 = _GEN_10622 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_16 = {_ans_17_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_18 = _ans_17_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_19 = _ans_17_leadingZeros_T_14 | _ans_17_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10623 = {{4'd0}, _ans_17_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_24 = _GEN_10623 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_26 = {_ans_17_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_28 = _ans_17_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_29 = _ans_17_leadingZeros_T_24 | _ans_17_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10624 = {{2'd0}, _ans_17_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_34 = _GEN_10624 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_36 = {_ans_17_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_38 = _ans_17_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_39 = _ans_17_leadingZeros_T_34 | _ans_17_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10625 = {{1'd0}, _ans_17_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_44 = _GEN_10625 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_46 = {_ans_17_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_48 = _ans_17_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_17_leadingZeros_T_49 = _ans_17_leadingZeros_T_44 | _ans_17_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10626 = {{8'd0}, ans_17_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_55 = _GEN_10626 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_57 = {ans_17_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_59 = _ans_17_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_60 = _ans_17_leadingZeros_T_55 | _ans_17_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10627 = {{4'd0}, _ans_17_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_65 = _GEN_10627 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_67 = {_ans_17_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_69 = _ans_17_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_70 = _ans_17_leadingZeros_T_65 | _ans_17_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10628 = {{2'd0}, _ans_17_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_75 = _GEN_10628 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_77 = {_ans_17_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_79 = _ans_17_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_80 = _ans_17_leadingZeros_T_75 | _ans_17_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10629 = {{1'd0}, _ans_17_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_85 = _GEN_10629 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_87 = {_ans_17_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_89 = _ans_17_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_17_leadingZeros_T_90 = _ans_17_leadingZeros_T_85 | _ans_17_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_17_leadingZeros_T_93 = {_ans_17_leadingZeros_T_49,_ans_17_leadingZeros_T_90,ans_17_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_17_leadingZeros_T_143 = _ans_17_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_144 = _ans_17_leadingZeros_T_93[46] ? 6'h2e : _ans_17_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_145 = _ans_17_leadingZeros_T_93[45] ? 6'h2d : _ans_17_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_146 = _ans_17_leadingZeros_T_93[44] ? 6'h2c : _ans_17_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_147 = _ans_17_leadingZeros_T_93[43] ? 6'h2b : _ans_17_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_148 = _ans_17_leadingZeros_T_93[42] ? 6'h2a : _ans_17_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_149 = _ans_17_leadingZeros_T_93[41] ? 6'h29 : _ans_17_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_150 = _ans_17_leadingZeros_T_93[40] ? 6'h28 : _ans_17_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_151 = _ans_17_leadingZeros_T_93[39] ? 6'h27 : _ans_17_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_152 = _ans_17_leadingZeros_T_93[38] ? 6'h26 : _ans_17_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_153 = _ans_17_leadingZeros_T_93[37] ? 6'h25 : _ans_17_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_154 = _ans_17_leadingZeros_T_93[36] ? 6'h24 : _ans_17_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_155 = _ans_17_leadingZeros_T_93[35] ? 6'h23 : _ans_17_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_156 = _ans_17_leadingZeros_T_93[34] ? 6'h22 : _ans_17_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_157 = _ans_17_leadingZeros_T_93[33] ? 6'h21 : _ans_17_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_158 = _ans_17_leadingZeros_T_93[32] ? 6'h20 : _ans_17_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_159 = _ans_17_leadingZeros_T_93[31] ? 6'h1f : _ans_17_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_160 = _ans_17_leadingZeros_T_93[30] ? 6'h1e : _ans_17_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_161 = _ans_17_leadingZeros_T_93[29] ? 6'h1d : _ans_17_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_162 = _ans_17_leadingZeros_T_93[28] ? 6'h1c : _ans_17_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_163 = _ans_17_leadingZeros_T_93[27] ? 6'h1b : _ans_17_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_164 = _ans_17_leadingZeros_T_93[26] ? 6'h1a : _ans_17_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_165 = _ans_17_leadingZeros_T_93[25] ? 6'h19 : _ans_17_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_166 = _ans_17_leadingZeros_T_93[24] ? 6'h18 : _ans_17_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_167 = _ans_17_leadingZeros_T_93[23] ? 6'h17 : _ans_17_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_168 = _ans_17_leadingZeros_T_93[22] ? 6'h16 : _ans_17_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_169 = _ans_17_leadingZeros_T_93[21] ? 6'h15 : _ans_17_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_170 = _ans_17_leadingZeros_T_93[20] ? 6'h14 : _ans_17_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_171 = _ans_17_leadingZeros_T_93[19] ? 6'h13 : _ans_17_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_172 = _ans_17_leadingZeros_T_93[18] ? 6'h12 : _ans_17_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_173 = _ans_17_leadingZeros_T_93[17] ? 6'h11 : _ans_17_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_174 = _ans_17_leadingZeros_T_93[16] ? 6'h10 : _ans_17_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_175 = _ans_17_leadingZeros_T_93[15] ? 6'hf : _ans_17_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_176 = _ans_17_leadingZeros_T_93[14] ? 6'he : _ans_17_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_177 = _ans_17_leadingZeros_T_93[13] ? 6'hd : _ans_17_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_178 = _ans_17_leadingZeros_T_93[12] ? 6'hc : _ans_17_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_179 = _ans_17_leadingZeros_T_93[11] ? 6'hb : _ans_17_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_180 = _ans_17_leadingZeros_T_93[10] ? 6'ha : _ans_17_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_181 = _ans_17_leadingZeros_T_93[9] ? 6'h9 : _ans_17_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_182 = _ans_17_leadingZeros_T_93[8] ? 6'h8 : _ans_17_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_183 = _ans_17_leadingZeros_T_93[7] ? 6'h7 : _ans_17_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_184 = _ans_17_leadingZeros_T_93[6] ? 6'h6 : _ans_17_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_185 = _ans_17_leadingZeros_T_93[5] ? 6'h5 : _ans_17_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_186 = _ans_17_leadingZeros_T_93[4] ? 6'h4 : _ans_17_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_187 = _ans_17_leadingZeros_T_93[3] ? 6'h3 : _ans_17_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_188 = _ans_17_leadingZeros_T_93[2] ? 6'h2 : _ans_17_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_189 = _ans_17_leadingZeros_T_93[1] ? 6'h1 : _ans_17_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_17_leadingZeros = _ans_17_leadingZeros_T_93[0] ? 6'h0 : _ans_17_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_expRaw_T_1 = 6'h1f - ans_17_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_17_expRaw = ans_17_isZero ? 6'h0 : _ans_17_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_17_shiftAmt_T_2 = ans_17_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_17_shiftAmt = ans_17_expRaw > 6'h3 ? _ans_17_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_17_mantissaRaw_T = ans_17_absClipped >> ans_17_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_17_mantissaRaw = _ans_17_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_17_mantissa = ans_17_expRaw >= 6'h3 ? ans_17_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_17_expAdjusted = ans_17_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_17_exp_T_4 = ans_17_expAdjusted > 7'hf ? 4'hf : ans_17_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_17_exp = ans_17_isZero ? 4'h0 : _ans_17_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_17_fp8 = {ans_17_clippedX[31],ans_17_exp,ans_17_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_18 = {24'h0,linear_bias_18}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_18 = tempSum_18 + biasExtended_18; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_18_sign = sum32_18[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_18_absX_T = ~sum32_18; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_18_absX_T_2 = _ans_18_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_18_absX = ans_18_sign ? _ans_18_absX_T_2 : sum32_18; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_18_shiftedX_T_1 = _GEN_10432 - ans_18_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_18_shiftedX_T_3 = ans_18_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_18_shiftedX = ans_18_sign ? _ans_18_shiftedX_T_1 : _ans_18_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_18_scaledX_T_1 = ans_18_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_18_scaledX = _ans_18_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_18_clippedX_T_2 = ans_18_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_18_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_18_clippedX = ans_18_scaledX > 49'h1c0 ? 49'h1c0 : _ans_18_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_18_absClipped_T_1 = ~ans_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_18_absClipped_T_3 = _ans_18_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_18_absClipped = ans_18_clippedX[31] ? _ans_18_absClipped_T_3 : ans_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_18_isZero = ans_18_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10632 = {{16'd0}, ans_18_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_4 = _GEN_10632 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_6 = {ans_18_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_8 = _ans_18_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_9 = _ans_18_leadingZeros_T_4 | _ans_18_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10633 = {{8'd0}, _ans_18_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_14 = _GEN_10633 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_16 = {_ans_18_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_18 = _ans_18_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_19 = _ans_18_leadingZeros_T_14 | _ans_18_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10634 = {{4'd0}, _ans_18_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_24 = _GEN_10634 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_26 = {_ans_18_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_28 = _ans_18_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_29 = _ans_18_leadingZeros_T_24 | _ans_18_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10635 = {{2'd0}, _ans_18_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_34 = _GEN_10635 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_36 = {_ans_18_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_38 = _ans_18_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_39 = _ans_18_leadingZeros_T_34 | _ans_18_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10636 = {{1'd0}, _ans_18_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_44 = _GEN_10636 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_46 = {_ans_18_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_48 = _ans_18_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_18_leadingZeros_T_49 = _ans_18_leadingZeros_T_44 | _ans_18_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10637 = {{8'd0}, ans_18_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_55 = _GEN_10637 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_57 = {ans_18_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_59 = _ans_18_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_60 = _ans_18_leadingZeros_T_55 | _ans_18_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10638 = {{4'd0}, _ans_18_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_65 = _GEN_10638 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_67 = {_ans_18_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_69 = _ans_18_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_70 = _ans_18_leadingZeros_T_65 | _ans_18_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10639 = {{2'd0}, _ans_18_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_75 = _GEN_10639 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_77 = {_ans_18_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_79 = _ans_18_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_80 = _ans_18_leadingZeros_T_75 | _ans_18_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10640 = {{1'd0}, _ans_18_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_85 = _GEN_10640 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_87 = {_ans_18_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_89 = _ans_18_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_18_leadingZeros_T_90 = _ans_18_leadingZeros_T_85 | _ans_18_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_18_leadingZeros_T_93 = {_ans_18_leadingZeros_T_49,_ans_18_leadingZeros_T_90,ans_18_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_18_leadingZeros_T_143 = _ans_18_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_144 = _ans_18_leadingZeros_T_93[46] ? 6'h2e : _ans_18_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_145 = _ans_18_leadingZeros_T_93[45] ? 6'h2d : _ans_18_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_146 = _ans_18_leadingZeros_T_93[44] ? 6'h2c : _ans_18_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_147 = _ans_18_leadingZeros_T_93[43] ? 6'h2b : _ans_18_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_148 = _ans_18_leadingZeros_T_93[42] ? 6'h2a : _ans_18_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_149 = _ans_18_leadingZeros_T_93[41] ? 6'h29 : _ans_18_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_150 = _ans_18_leadingZeros_T_93[40] ? 6'h28 : _ans_18_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_151 = _ans_18_leadingZeros_T_93[39] ? 6'h27 : _ans_18_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_152 = _ans_18_leadingZeros_T_93[38] ? 6'h26 : _ans_18_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_153 = _ans_18_leadingZeros_T_93[37] ? 6'h25 : _ans_18_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_154 = _ans_18_leadingZeros_T_93[36] ? 6'h24 : _ans_18_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_155 = _ans_18_leadingZeros_T_93[35] ? 6'h23 : _ans_18_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_156 = _ans_18_leadingZeros_T_93[34] ? 6'h22 : _ans_18_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_157 = _ans_18_leadingZeros_T_93[33] ? 6'h21 : _ans_18_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_158 = _ans_18_leadingZeros_T_93[32] ? 6'h20 : _ans_18_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_159 = _ans_18_leadingZeros_T_93[31] ? 6'h1f : _ans_18_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_160 = _ans_18_leadingZeros_T_93[30] ? 6'h1e : _ans_18_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_161 = _ans_18_leadingZeros_T_93[29] ? 6'h1d : _ans_18_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_162 = _ans_18_leadingZeros_T_93[28] ? 6'h1c : _ans_18_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_163 = _ans_18_leadingZeros_T_93[27] ? 6'h1b : _ans_18_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_164 = _ans_18_leadingZeros_T_93[26] ? 6'h1a : _ans_18_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_165 = _ans_18_leadingZeros_T_93[25] ? 6'h19 : _ans_18_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_166 = _ans_18_leadingZeros_T_93[24] ? 6'h18 : _ans_18_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_167 = _ans_18_leadingZeros_T_93[23] ? 6'h17 : _ans_18_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_168 = _ans_18_leadingZeros_T_93[22] ? 6'h16 : _ans_18_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_169 = _ans_18_leadingZeros_T_93[21] ? 6'h15 : _ans_18_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_170 = _ans_18_leadingZeros_T_93[20] ? 6'h14 : _ans_18_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_171 = _ans_18_leadingZeros_T_93[19] ? 6'h13 : _ans_18_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_172 = _ans_18_leadingZeros_T_93[18] ? 6'h12 : _ans_18_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_173 = _ans_18_leadingZeros_T_93[17] ? 6'h11 : _ans_18_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_174 = _ans_18_leadingZeros_T_93[16] ? 6'h10 : _ans_18_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_175 = _ans_18_leadingZeros_T_93[15] ? 6'hf : _ans_18_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_176 = _ans_18_leadingZeros_T_93[14] ? 6'he : _ans_18_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_177 = _ans_18_leadingZeros_T_93[13] ? 6'hd : _ans_18_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_178 = _ans_18_leadingZeros_T_93[12] ? 6'hc : _ans_18_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_179 = _ans_18_leadingZeros_T_93[11] ? 6'hb : _ans_18_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_180 = _ans_18_leadingZeros_T_93[10] ? 6'ha : _ans_18_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_181 = _ans_18_leadingZeros_T_93[9] ? 6'h9 : _ans_18_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_182 = _ans_18_leadingZeros_T_93[8] ? 6'h8 : _ans_18_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_183 = _ans_18_leadingZeros_T_93[7] ? 6'h7 : _ans_18_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_184 = _ans_18_leadingZeros_T_93[6] ? 6'h6 : _ans_18_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_185 = _ans_18_leadingZeros_T_93[5] ? 6'h5 : _ans_18_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_186 = _ans_18_leadingZeros_T_93[4] ? 6'h4 : _ans_18_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_187 = _ans_18_leadingZeros_T_93[3] ? 6'h3 : _ans_18_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_188 = _ans_18_leadingZeros_T_93[2] ? 6'h2 : _ans_18_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_189 = _ans_18_leadingZeros_T_93[1] ? 6'h1 : _ans_18_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_18_leadingZeros = _ans_18_leadingZeros_T_93[0] ? 6'h0 : _ans_18_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_expRaw_T_1 = 6'h1f - ans_18_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_18_expRaw = ans_18_isZero ? 6'h0 : _ans_18_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_18_shiftAmt_T_2 = ans_18_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_18_shiftAmt = ans_18_expRaw > 6'h3 ? _ans_18_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_18_mantissaRaw_T = ans_18_absClipped >> ans_18_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_18_mantissaRaw = _ans_18_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_18_mantissa = ans_18_expRaw >= 6'h3 ? ans_18_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_18_expAdjusted = ans_18_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_18_exp_T_4 = ans_18_expAdjusted > 7'hf ? 4'hf : ans_18_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_18_exp = ans_18_isZero ? 4'h0 : _ans_18_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_18_fp8 = {ans_18_clippedX[31],ans_18_exp,ans_18_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_19 = {24'h0,linear_bias_19}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_19 = tempSum_19 + biasExtended_19; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_19_sign = sum32_19[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_19_absX_T = ~sum32_19; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_19_absX_T_2 = _ans_19_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_19_absX = ans_19_sign ? _ans_19_absX_T_2 : sum32_19; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_19_shiftedX_T_1 = _GEN_10432 - ans_19_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_19_shiftedX_T_3 = ans_19_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_19_shiftedX = ans_19_sign ? _ans_19_shiftedX_T_1 : _ans_19_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_19_scaledX_T_1 = ans_19_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_19_scaledX = _ans_19_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_19_clippedX_T_2 = ans_19_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_19_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_19_clippedX = ans_19_scaledX > 49'h1c0 ? 49'h1c0 : _ans_19_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_19_absClipped_T_1 = ~ans_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_19_absClipped_T_3 = _ans_19_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_19_absClipped = ans_19_clippedX[31] ? _ans_19_absClipped_T_3 : ans_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_19_isZero = ans_19_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10643 = {{16'd0}, ans_19_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_4 = _GEN_10643 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_6 = {ans_19_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_8 = _ans_19_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_9 = _ans_19_leadingZeros_T_4 | _ans_19_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10644 = {{8'd0}, _ans_19_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_14 = _GEN_10644 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_16 = {_ans_19_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_18 = _ans_19_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_19 = _ans_19_leadingZeros_T_14 | _ans_19_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10645 = {{4'd0}, _ans_19_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_24 = _GEN_10645 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_26 = {_ans_19_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_28 = _ans_19_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_29 = _ans_19_leadingZeros_T_24 | _ans_19_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10646 = {{2'd0}, _ans_19_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_34 = _GEN_10646 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_36 = {_ans_19_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_38 = _ans_19_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_39 = _ans_19_leadingZeros_T_34 | _ans_19_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10647 = {{1'd0}, _ans_19_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_44 = _GEN_10647 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_46 = {_ans_19_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_48 = _ans_19_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_19_leadingZeros_T_49 = _ans_19_leadingZeros_T_44 | _ans_19_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10648 = {{8'd0}, ans_19_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_55 = _GEN_10648 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_57 = {ans_19_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_59 = _ans_19_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_60 = _ans_19_leadingZeros_T_55 | _ans_19_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10649 = {{4'd0}, _ans_19_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_65 = _GEN_10649 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_67 = {_ans_19_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_69 = _ans_19_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_70 = _ans_19_leadingZeros_T_65 | _ans_19_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10650 = {{2'd0}, _ans_19_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_75 = _GEN_10650 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_77 = {_ans_19_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_79 = _ans_19_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_80 = _ans_19_leadingZeros_T_75 | _ans_19_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10651 = {{1'd0}, _ans_19_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_85 = _GEN_10651 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_87 = {_ans_19_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_89 = _ans_19_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_19_leadingZeros_T_90 = _ans_19_leadingZeros_T_85 | _ans_19_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_19_leadingZeros_T_93 = {_ans_19_leadingZeros_T_49,_ans_19_leadingZeros_T_90,ans_19_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_19_leadingZeros_T_143 = _ans_19_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_144 = _ans_19_leadingZeros_T_93[46] ? 6'h2e : _ans_19_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_145 = _ans_19_leadingZeros_T_93[45] ? 6'h2d : _ans_19_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_146 = _ans_19_leadingZeros_T_93[44] ? 6'h2c : _ans_19_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_147 = _ans_19_leadingZeros_T_93[43] ? 6'h2b : _ans_19_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_148 = _ans_19_leadingZeros_T_93[42] ? 6'h2a : _ans_19_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_149 = _ans_19_leadingZeros_T_93[41] ? 6'h29 : _ans_19_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_150 = _ans_19_leadingZeros_T_93[40] ? 6'h28 : _ans_19_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_151 = _ans_19_leadingZeros_T_93[39] ? 6'h27 : _ans_19_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_152 = _ans_19_leadingZeros_T_93[38] ? 6'h26 : _ans_19_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_153 = _ans_19_leadingZeros_T_93[37] ? 6'h25 : _ans_19_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_154 = _ans_19_leadingZeros_T_93[36] ? 6'h24 : _ans_19_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_155 = _ans_19_leadingZeros_T_93[35] ? 6'h23 : _ans_19_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_156 = _ans_19_leadingZeros_T_93[34] ? 6'h22 : _ans_19_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_157 = _ans_19_leadingZeros_T_93[33] ? 6'h21 : _ans_19_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_158 = _ans_19_leadingZeros_T_93[32] ? 6'h20 : _ans_19_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_159 = _ans_19_leadingZeros_T_93[31] ? 6'h1f : _ans_19_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_160 = _ans_19_leadingZeros_T_93[30] ? 6'h1e : _ans_19_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_161 = _ans_19_leadingZeros_T_93[29] ? 6'h1d : _ans_19_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_162 = _ans_19_leadingZeros_T_93[28] ? 6'h1c : _ans_19_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_163 = _ans_19_leadingZeros_T_93[27] ? 6'h1b : _ans_19_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_164 = _ans_19_leadingZeros_T_93[26] ? 6'h1a : _ans_19_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_165 = _ans_19_leadingZeros_T_93[25] ? 6'h19 : _ans_19_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_166 = _ans_19_leadingZeros_T_93[24] ? 6'h18 : _ans_19_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_167 = _ans_19_leadingZeros_T_93[23] ? 6'h17 : _ans_19_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_168 = _ans_19_leadingZeros_T_93[22] ? 6'h16 : _ans_19_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_169 = _ans_19_leadingZeros_T_93[21] ? 6'h15 : _ans_19_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_170 = _ans_19_leadingZeros_T_93[20] ? 6'h14 : _ans_19_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_171 = _ans_19_leadingZeros_T_93[19] ? 6'h13 : _ans_19_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_172 = _ans_19_leadingZeros_T_93[18] ? 6'h12 : _ans_19_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_173 = _ans_19_leadingZeros_T_93[17] ? 6'h11 : _ans_19_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_174 = _ans_19_leadingZeros_T_93[16] ? 6'h10 : _ans_19_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_175 = _ans_19_leadingZeros_T_93[15] ? 6'hf : _ans_19_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_176 = _ans_19_leadingZeros_T_93[14] ? 6'he : _ans_19_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_177 = _ans_19_leadingZeros_T_93[13] ? 6'hd : _ans_19_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_178 = _ans_19_leadingZeros_T_93[12] ? 6'hc : _ans_19_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_179 = _ans_19_leadingZeros_T_93[11] ? 6'hb : _ans_19_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_180 = _ans_19_leadingZeros_T_93[10] ? 6'ha : _ans_19_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_181 = _ans_19_leadingZeros_T_93[9] ? 6'h9 : _ans_19_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_182 = _ans_19_leadingZeros_T_93[8] ? 6'h8 : _ans_19_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_183 = _ans_19_leadingZeros_T_93[7] ? 6'h7 : _ans_19_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_184 = _ans_19_leadingZeros_T_93[6] ? 6'h6 : _ans_19_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_185 = _ans_19_leadingZeros_T_93[5] ? 6'h5 : _ans_19_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_186 = _ans_19_leadingZeros_T_93[4] ? 6'h4 : _ans_19_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_187 = _ans_19_leadingZeros_T_93[3] ? 6'h3 : _ans_19_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_188 = _ans_19_leadingZeros_T_93[2] ? 6'h2 : _ans_19_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_189 = _ans_19_leadingZeros_T_93[1] ? 6'h1 : _ans_19_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_19_leadingZeros = _ans_19_leadingZeros_T_93[0] ? 6'h0 : _ans_19_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_expRaw_T_1 = 6'h1f - ans_19_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_19_expRaw = ans_19_isZero ? 6'h0 : _ans_19_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_19_shiftAmt_T_2 = ans_19_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_19_shiftAmt = ans_19_expRaw > 6'h3 ? _ans_19_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_19_mantissaRaw_T = ans_19_absClipped >> ans_19_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_19_mantissaRaw = _ans_19_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_19_mantissa = ans_19_expRaw >= 6'h3 ? ans_19_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_19_expAdjusted = ans_19_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_19_exp_T_4 = ans_19_expAdjusted > 7'hf ? 4'hf : ans_19_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_19_exp = ans_19_isZero ? 4'h0 : _ans_19_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_19_fp8 = {ans_19_clippedX[31],ans_19_exp,ans_19_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_20 = {24'h0,linear_bias_20}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_20 = tempSum_20 + biasExtended_20; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_20_sign = sum32_20[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_20_absX_T = ~sum32_20; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_20_absX_T_2 = _ans_20_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_20_absX = ans_20_sign ? _ans_20_absX_T_2 : sum32_20; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_20_shiftedX_T_1 = _GEN_10432 - ans_20_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_20_shiftedX_T_3 = ans_20_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_20_shiftedX = ans_20_sign ? _ans_20_shiftedX_T_1 : _ans_20_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_20_scaledX_T_1 = ans_20_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_20_scaledX = _ans_20_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_20_clippedX_T_2 = ans_20_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_20_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_20_clippedX = ans_20_scaledX > 49'h1c0 ? 49'h1c0 : _ans_20_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_20_absClipped_T_1 = ~ans_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_20_absClipped_T_3 = _ans_20_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_20_absClipped = ans_20_clippedX[31] ? _ans_20_absClipped_T_3 : ans_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_20_isZero = ans_20_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10654 = {{16'd0}, ans_20_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_4 = _GEN_10654 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_6 = {ans_20_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_8 = _ans_20_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_9 = _ans_20_leadingZeros_T_4 | _ans_20_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10655 = {{8'd0}, _ans_20_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_14 = _GEN_10655 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_16 = {_ans_20_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_18 = _ans_20_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_19 = _ans_20_leadingZeros_T_14 | _ans_20_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10656 = {{4'd0}, _ans_20_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_24 = _GEN_10656 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_26 = {_ans_20_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_28 = _ans_20_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_29 = _ans_20_leadingZeros_T_24 | _ans_20_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10657 = {{2'd0}, _ans_20_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_34 = _GEN_10657 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_36 = {_ans_20_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_38 = _ans_20_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_39 = _ans_20_leadingZeros_T_34 | _ans_20_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10658 = {{1'd0}, _ans_20_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_44 = _GEN_10658 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_46 = {_ans_20_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_48 = _ans_20_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_20_leadingZeros_T_49 = _ans_20_leadingZeros_T_44 | _ans_20_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10659 = {{8'd0}, ans_20_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_55 = _GEN_10659 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_57 = {ans_20_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_59 = _ans_20_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_60 = _ans_20_leadingZeros_T_55 | _ans_20_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10660 = {{4'd0}, _ans_20_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_65 = _GEN_10660 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_67 = {_ans_20_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_69 = _ans_20_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_70 = _ans_20_leadingZeros_T_65 | _ans_20_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10661 = {{2'd0}, _ans_20_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_75 = _GEN_10661 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_77 = {_ans_20_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_79 = _ans_20_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_80 = _ans_20_leadingZeros_T_75 | _ans_20_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10662 = {{1'd0}, _ans_20_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_85 = _GEN_10662 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_87 = {_ans_20_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_89 = _ans_20_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_20_leadingZeros_T_90 = _ans_20_leadingZeros_T_85 | _ans_20_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_20_leadingZeros_T_93 = {_ans_20_leadingZeros_T_49,_ans_20_leadingZeros_T_90,ans_20_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_20_leadingZeros_T_143 = _ans_20_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_144 = _ans_20_leadingZeros_T_93[46] ? 6'h2e : _ans_20_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_145 = _ans_20_leadingZeros_T_93[45] ? 6'h2d : _ans_20_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_146 = _ans_20_leadingZeros_T_93[44] ? 6'h2c : _ans_20_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_147 = _ans_20_leadingZeros_T_93[43] ? 6'h2b : _ans_20_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_148 = _ans_20_leadingZeros_T_93[42] ? 6'h2a : _ans_20_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_149 = _ans_20_leadingZeros_T_93[41] ? 6'h29 : _ans_20_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_150 = _ans_20_leadingZeros_T_93[40] ? 6'h28 : _ans_20_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_151 = _ans_20_leadingZeros_T_93[39] ? 6'h27 : _ans_20_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_152 = _ans_20_leadingZeros_T_93[38] ? 6'h26 : _ans_20_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_153 = _ans_20_leadingZeros_T_93[37] ? 6'h25 : _ans_20_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_154 = _ans_20_leadingZeros_T_93[36] ? 6'h24 : _ans_20_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_155 = _ans_20_leadingZeros_T_93[35] ? 6'h23 : _ans_20_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_156 = _ans_20_leadingZeros_T_93[34] ? 6'h22 : _ans_20_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_157 = _ans_20_leadingZeros_T_93[33] ? 6'h21 : _ans_20_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_158 = _ans_20_leadingZeros_T_93[32] ? 6'h20 : _ans_20_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_159 = _ans_20_leadingZeros_T_93[31] ? 6'h1f : _ans_20_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_160 = _ans_20_leadingZeros_T_93[30] ? 6'h1e : _ans_20_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_161 = _ans_20_leadingZeros_T_93[29] ? 6'h1d : _ans_20_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_162 = _ans_20_leadingZeros_T_93[28] ? 6'h1c : _ans_20_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_163 = _ans_20_leadingZeros_T_93[27] ? 6'h1b : _ans_20_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_164 = _ans_20_leadingZeros_T_93[26] ? 6'h1a : _ans_20_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_165 = _ans_20_leadingZeros_T_93[25] ? 6'h19 : _ans_20_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_166 = _ans_20_leadingZeros_T_93[24] ? 6'h18 : _ans_20_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_167 = _ans_20_leadingZeros_T_93[23] ? 6'h17 : _ans_20_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_168 = _ans_20_leadingZeros_T_93[22] ? 6'h16 : _ans_20_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_169 = _ans_20_leadingZeros_T_93[21] ? 6'h15 : _ans_20_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_170 = _ans_20_leadingZeros_T_93[20] ? 6'h14 : _ans_20_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_171 = _ans_20_leadingZeros_T_93[19] ? 6'h13 : _ans_20_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_172 = _ans_20_leadingZeros_T_93[18] ? 6'h12 : _ans_20_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_173 = _ans_20_leadingZeros_T_93[17] ? 6'h11 : _ans_20_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_174 = _ans_20_leadingZeros_T_93[16] ? 6'h10 : _ans_20_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_175 = _ans_20_leadingZeros_T_93[15] ? 6'hf : _ans_20_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_176 = _ans_20_leadingZeros_T_93[14] ? 6'he : _ans_20_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_177 = _ans_20_leadingZeros_T_93[13] ? 6'hd : _ans_20_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_178 = _ans_20_leadingZeros_T_93[12] ? 6'hc : _ans_20_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_179 = _ans_20_leadingZeros_T_93[11] ? 6'hb : _ans_20_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_180 = _ans_20_leadingZeros_T_93[10] ? 6'ha : _ans_20_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_181 = _ans_20_leadingZeros_T_93[9] ? 6'h9 : _ans_20_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_182 = _ans_20_leadingZeros_T_93[8] ? 6'h8 : _ans_20_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_183 = _ans_20_leadingZeros_T_93[7] ? 6'h7 : _ans_20_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_184 = _ans_20_leadingZeros_T_93[6] ? 6'h6 : _ans_20_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_185 = _ans_20_leadingZeros_T_93[5] ? 6'h5 : _ans_20_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_186 = _ans_20_leadingZeros_T_93[4] ? 6'h4 : _ans_20_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_187 = _ans_20_leadingZeros_T_93[3] ? 6'h3 : _ans_20_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_188 = _ans_20_leadingZeros_T_93[2] ? 6'h2 : _ans_20_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_189 = _ans_20_leadingZeros_T_93[1] ? 6'h1 : _ans_20_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_20_leadingZeros = _ans_20_leadingZeros_T_93[0] ? 6'h0 : _ans_20_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_expRaw_T_1 = 6'h1f - ans_20_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_20_expRaw = ans_20_isZero ? 6'h0 : _ans_20_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_20_shiftAmt_T_2 = ans_20_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_20_shiftAmt = ans_20_expRaw > 6'h3 ? _ans_20_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_20_mantissaRaw_T = ans_20_absClipped >> ans_20_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_20_mantissaRaw = _ans_20_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_20_mantissa = ans_20_expRaw >= 6'h3 ? ans_20_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_20_expAdjusted = ans_20_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_20_exp_T_4 = ans_20_expAdjusted > 7'hf ? 4'hf : ans_20_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_20_exp = ans_20_isZero ? 4'h0 : _ans_20_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_20_fp8 = {ans_20_clippedX[31],ans_20_exp,ans_20_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_21 = {24'h0,linear_bias_21}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_21 = tempSum_21 + biasExtended_21; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_21_sign = sum32_21[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_21_absX_T = ~sum32_21; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_21_absX_T_2 = _ans_21_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_21_absX = ans_21_sign ? _ans_21_absX_T_2 : sum32_21; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_21_shiftedX_T_1 = _GEN_10432 - ans_21_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_21_shiftedX_T_3 = ans_21_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_21_shiftedX = ans_21_sign ? _ans_21_shiftedX_T_1 : _ans_21_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_21_scaledX_T_1 = ans_21_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_21_scaledX = _ans_21_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_21_clippedX_T_2 = ans_21_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_21_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_21_clippedX = ans_21_scaledX > 49'h1c0 ? 49'h1c0 : _ans_21_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_21_absClipped_T_1 = ~ans_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_21_absClipped_T_3 = _ans_21_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_21_absClipped = ans_21_clippedX[31] ? _ans_21_absClipped_T_3 : ans_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_21_isZero = ans_21_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10665 = {{16'd0}, ans_21_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_4 = _GEN_10665 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_6 = {ans_21_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_8 = _ans_21_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_9 = _ans_21_leadingZeros_T_4 | _ans_21_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10666 = {{8'd0}, _ans_21_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_14 = _GEN_10666 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_16 = {_ans_21_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_18 = _ans_21_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_19 = _ans_21_leadingZeros_T_14 | _ans_21_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10667 = {{4'd0}, _ans_21_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_24 = _GEN_10667 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_26 = {_ans_21_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_28 = _ans_21_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_29 = _ans_21_leadingZeros_T_24 | _ans_21_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10668 = {{2'd0}, _ans_21_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_34 = _GEN_10668 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_36 = {_ans_21_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_38 = _ans_21_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_39 = _ans_21_leadingZeros_T_34 | _ans_21_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10669 = {{1'd0}, _ans_21_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_44 = _GEN_10669 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_46 = {_ans_21_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_48 = _ans_21_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_21_leadingZeros_T_49 = _ans_21_leadingZeros_T_44 | _ans_21_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10670 = {{8'd0}, ans_21_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_55 = _GEN_10670 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_57 = {ans_21_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_59 = _ans_21_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_60 = _ans_21_leadingZeros_T_55 | _ans_21_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10671 = {{4'd0}, _ans_21_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_65 = _GEN_10671 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_67 = {_ans_21_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_69 = _ans_21_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_70 = _ans_21_leadingZeros_T_65 | _ans_21_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10672 = {{2'd0}, _ans_21_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_75 = _GEN_10672 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_77 = {_ans_21_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_79 = _ans_21_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_80 = _ans_21_leadingZeros_T_75 | _ans_21_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10673 = {{1'd0}, _ans_21_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_85 = _GEN_10673 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_87 = {_ans_21_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_89 = _ans_21_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_21_leadingZeros_T_90 = _ans_21_leadingZeros_T_85 | _ans_21_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_21_leadingZeros_T_93 = {_ans_21_leadingZeros_T_49,_ans_21_leadingZeros_T_90,ans_21_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_21_leadingZeros_T_143 = _ans_21_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_144 = _ans_21_leadingZeros_T_93[46] ? 6'h2e : _ans_21_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_145 = _ans_21_leadingZeros_T_93[45] ? 6'h2d : _ans_21_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_146 = _ans_21_leadingZeros_T_93[44] ? 6'h2c : _ans_21_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_147 = _ans_21_leadingZeros_T_93[43] ? 6'h2b : _ans_21_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_148 = _ans_21_leadingZeros_T_93[42] ? 6'h2a : _ans_21_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_149 = _ans_21_leadingZeros_T_93[41] ? 6'h29 : _ans_21_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_150 = _ans_21_leadingZeros_T_93[40] ? 6'h28 : _ans_21_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_151 = _ans_21_leadingZeros_T_93[39] ? 6'h27 : _ans_21_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_152 = _ans_21_leadingZeros_T_93[38] ? 6'h26 : _ans_21_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_153 = _ans_21_leadingZeros_T_93[37] ? 6'h25 : _ans_21_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_154 = _ans_21_leadingZeros_T_93[36] ? 6'h24 : _ans_21_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_155 = _ans_21_leadingZeros_T_93[35] ? 6'h23 : _ans_21_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_156 = _ans_21_leadingZeros_T_93[34] ? 6'h22 : _ans_21_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_157 = _ans_21_leadingZeros_T_93[33] ? 6'h21 : _ans_21_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_158 = _ans_21_leadingZeros_T_93[32] ? 6'h20 : _ans_21_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_159 = _ans_21_leadingZeros_T_93[31] ? 6'h1f : _ans_21_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_160 = _ans_21_leadingZeros_T_93[30] ? 6'h1e : _ans_21_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_161 = _ans_21_leadingZeros_T_93[29] ? 6'h1d : _ans_21_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_162 = _ans_21_leadingZeros_T_93[28] ? 6'h1c : _ans_21_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_163 = _ans_21_leadingZeros_T_93[27] ? 6'h1b : _ans_21_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_164 = _ans_21_leadingZeros_T_93[26] ? 6'h1a : _ans_21_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_165 = _ans_21_leadingZeros_T_93[25] ? 6'h19 : _ans_21_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_166 = _ans_21_leadingZeros_T_93[24] ? 6'h18 : _ans_21_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_167 = _ans_21_leadingZeros_T_93[23] ? 6'h17 : _ans_21_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_168 = _ans_21_leadingZeros_T_93[22] ? 6'h16 : _ans_21_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_169 = _ans_21_leadingZeros_T_93[21] ? 6'h15 : _ans_21_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_170 = _ans_21_leadingZeros_T_93[20] ? 6'h14 : _ans_21_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_171 = _ans_21_leadingZeros_T_93[19] ? 6'h13 : _ans_21_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_172 = _ans_21_leadingZeros_T_93[18] ? 6'h12 : _ans_21_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_173 = _ans_21_leadingZeros_T_93[17] ? 6'h11 : _ans_21_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_174 = _ans_21_leadingZeros_T_93[16] ? 6'h10 : _ans_21_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_175 = _ans_21_leadingZeros_T_93[15] ? 6'hf : _ans_21_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_176 = _ans_21_leadingZeros_T_93[14] ? 6'he : _ans_21_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_177 = _ans_21_leadingZeros_T_93[13] ? 6'hd : _ans_21_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_178 = _ans_21_leadingZeros_T_93[12] ? 6'hc : _ans_21_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_179 = _ans_21_leadingZeros_T_93[11] ? 6'hb : _ans_21_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_180 = _ans_21_leadingZeros_T_93[10] ? 6'ha : _ans_21_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_181 = _ans_21_leadingZeros_T_93[9] ? 6'h9 : _ans_21_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_182 = _ans_21_leadingZeros_T_93[8] ? 6'h8 : _ans_21_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_183 = _ans_21_leadingZeros_T_93[7] ? 6'h7 : _ans_21_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_184 = _ans_21_leadingZeros_T_93[6] ? 6'h6 : _ans_21_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_185 = _ans_21_leadingZeros_T_93[5] ? 6'h5 : _ans_21_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_186 = _ans_21_leadingZeros_T_93[4] ? 6'h4 : _ans_21_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_187 = _ans_21_leadingZeros_T_93[3] ? 6'h3 : _ans_21_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_188 = _ans_21_leadingZeros_T_93[2] ? 6'h2 : _ans_21_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_189 = _ans_21_leadingZeros_T_93[1] ? 6'h1 : _ans_21_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_21_leadingZeros = _ans_21_leadingZeros_T_93[0] ? 6'h0 : _ans_21_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_expRaw_T_1 = 6'h1f - ans_21_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_21_expRaw = ans_21_isZero ? 6'h0 : _ans_21_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_21_shiftAmt_T_2 = ans_21_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_21_shiftAmt = ans_21_expRaw > 6'h3 ? _ans_21_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_21_mantissaRaw_T = ans_21_absClipped >> ans_21_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_21_mantissaRaw = _ans_21_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_21_mantissa = ans_21_expRaw >= 6'h3 ? ans_21_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_21_expAdjusted = ans_21_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_21_exp_T_4 = ans_21_expAdjusted > 7'hf ? 4'hf : ans_21_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_21_exp = ans_21_isZero ? 4'h0 : _ans_21_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_21_fp8 = {ans_21_clippedX[31],ans_21_exp,ans_21_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_22 = {24'h0,linear_bias_22}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_22 = tempSum_22 + biasExtended_22; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_22_sign = sum32_22[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_22_absX_T = ~sum32_22; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_22_absX_T_2 = _ans_22_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_22_absX = ans_22_sign ? _ans_22_absX_T_2 : sum32_22; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_22_shiftedX_T_1 = _GEN_10432 - ans_22_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_22_shiftedX_T_3 = ans_22_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_22_shiftedX = ans_22_sign ? _ans_22_shiftedX_T_1 : _ans_22_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_22_scaledX_T_1 = ans_22_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_22_scaledX = _ans_22_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_22_clippedX_T_2 = ans_22_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_22_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_22_clippedX = ans_22_scaledX > 49'h1c0 ? 49'h1c0 : _ans_22_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_22_absClipped_T_1 = ~ans_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_22_absClipped_T_3 = _ans_22_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_22_absClipped = ans_22_clippedX[31] ? _ans_22_absClipped_T_3 : ans_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_22_isZero = ans_22_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10676 = {{16'd0}, ans_22_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_4 = _GEN_10676 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_6 = {ans_22_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_8 = _ans_22_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_9 = _ans_22_leadingZeros_T_4 | _ans_22_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10677 = {{8'd0}, _ans_22_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_14 = _GEN_10677 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_16 = {_ans_22_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_18 = _ans_22_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_19 = _ans_22_leadingZeros_T_14 | _ans_22_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10678 = {{4'd0}, _ans_22_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_24 = _GEN_10678 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_26 = {_ans_22_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_28 = _ans_22_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_29 = _ans_22_leadingZeros_T_24 | _ans_22_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10679 = {{2'd0}, _ans_22_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_34 = _GEN_10679 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_36 = {_ans_22_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_38 = _ans_22_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_39 = _ans_22_leadingZeros_T_34 | _ans_22_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10680 = {{1'd0}, _ans_22_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_44 = _GEN_10680 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_46 = {_ans_22_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_48 = _ans_22_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_22_leadingZeros_T_49 = _ans_22_leadingZeros_T_44 | _ans_22_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10681 = {{8'd0}, ans_22_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_55 = _GEN_10681 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_57 = {ans_22_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_59 = _ans_22_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_60 = _ans_22_leadingZeros_T_55 | _ans_22_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10682 = {{4'd0}, _ans_22_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_65 = _GEN_10682 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_67 = {_ans_22_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_69 = _ans_22_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_70 = _ans_22_leadingZeros_T_65 | _ans_22_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10683 = {{2'd0}, _ans_22_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_75 = _GEN_10683 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_77 = {_ans_22_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_79 = _ans_22_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_80 = _ans_22_leadingZeros_T_75 | _ans_22_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10684 = {{1'd0}, _ans_22_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_85 = _GEN_10684 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_87 = {_ans_22_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_89 = _ans_22_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_22_leadingZeros_T_90 = _ans_22_leadingZeros_T_85 | _ans_22_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_22_leadingZeros_T_93 = {_ans_22_leadingZeros_T_49,_ans_22_leadingZeros_T_90,ans_22_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_22_leadingZeros_T_143 = _ans_22_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_144 = _ans_22_leadingZeros_T_93[46] ? 6'h2e : _ans_22_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_145 = _ans_22_leadingZeros_T_93[45] ? 6'h2d : _ans_22_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_146 = _ans_22_leadingZeros_T_93[44] ? 6'h2c : _ans_22_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_147 = _ans_22_leadingZeros_T_93[43] ? 6'h2b : _ans_22_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_148 = _ans_22_leadingZeros_T_93[42] ? 6'h2a : _ans_22_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_149 = _ans_22_leadingZeros_T_93[41] ? 6'h29 : _ans_22_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_150 = _ans_22_leadingZeros_T_93[40] ? 6'h28 : _ans_22_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_151 = _ans_22_leadingZeros_T_93[39] ? 6'h27 : _ans_22_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_152 = _ans_22_leadingZeros_T_93[38] ? 6'h26 : _ans_22_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_153 = _ans_22_leadingZeros_T_93[37] ? 6'h25 : _ans_22_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_154 = _ans_22_leadingZeros_T_93[36] ? 6'h24 : _ans_22_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_155 = _ans_22_leadingZeros_T_93[35] ? 6'h23 : _ans_22_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_156 = _ans_22_leadingZeros_T_93[34] ? 6'h22 : _ans_22_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_157 = _ans_22_leadingZeros_T_93[33] ? 6'h21 : _ans_22_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_158 = _ans_22_leadingZeros_T_93[32] ? 6'h20 : _ans_22_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_159 = _ans_22_leadingZeros_T_93[31] ? 6'h1f : _ans_22_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_160 = _ans_22_leadingZeros_T_93[30] ? 6'h1e : _ans_22_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_161 = _ans_22_leadingZeros_T_93[29] ? 6'h1d : _ans_22_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_162 = _ans_22_leadingZeros_T_93[28] ? 6'h1c : _ans_22_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_163 = _ans_22_leadingZeros_T_93[27] ? 6'h1b : _ans_22_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_164 = _ans_22_leadingZeros_T_93[26] ? 6'h1a : _ans_22_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_165 = _ans_22_leadingZeros_T_93[25] ? 6'h19 : _ans_22_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_166 = _ans_22_leadingZeros_T_93[24] ? 6'h18 : _ans_22_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_167 = _ans_22_leadingZeros_T_93[23] ? 6'h17 : _ans_22_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_168 = _ans_22_leadingZeros_T_93[22] ? 6'h16 : _ans_22_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_169 = _ans_22_leadingZeros_T_93[21] ? 6'h15 : _ans_22_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_170 = _ans_22_leadingZeros_T_93[20] ? 6'h14 : _ans_22_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_171 = _ans_22_leadingZeros_T_93[19] ? 6'h13 : _ans_22_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_172 = _ans_22_leadingZeros_T_93[18] ? 6'h12 : _ans_22_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_173 = _ans_22_leadingZeros_T_93[17] ? 6'h11 : _ans_22_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_174 = _ans_22_leadingZeros_T_93[16] ? 6'h10 : _ans_22_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_175 = _ans_22_leadingZeros_T_93[15] ? 6'hf : _ans_22_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_176 = _ans_22_leadingZeros_T_93[14] ? 6'he : _ans_22_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_177 = _ans_22_leadingZeros_T_93[13] ? 6'hd : _ans_22_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_178 = _ans_22_leadingZeros_T_93[12] ? 6'hc : _ans_22_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_179 = _ans_22_leadingZeros_T_93[11] ? 6'hb : _ans_22_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_180 = _ans_22_leadingZeros_T_93[10] ? 6'ha : _ans_22_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_181 = _ans_22_leadingZeros_T_93[9] ? 6'h9 : _ans_22_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_182 = _ans_22_leadingZeros_T_93[8] ? 6'h8 : _ans_22_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_183 = _ans_22_leadingZeros_T_93[7] ? 6'h7 : _ans_22_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_184 = _ans_22_leadingZeros_T_93[6] ? 6'h6 : _ans_22_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_185 = _ans_22_leadingZeros_T_93[5] ? 6'h5 : _ans_22_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_186 = _ans_22_leadingZeros_T_93[4] ? 6'h4 : _ans_22_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_187 = _ans_22_leadingZeros_T_93[3] ? 6'h3 : _ans_22_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_188 = _ans_22_leadingZeros_T_93[2] ? 6'h2 : _ans_22_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_189 = _ans_22_leadingZeros_T_93[1] ? 6'h1 : _ans_22_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_22_leadingZeros = _ans_22_leadingZeros_T_93[0] ? 6'h0 : _ans_22_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_expRaw_T_1 = 6'h1f - ans_22_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_22_expRaw = ans_22_isZero ? 6'h0 : _ans_22_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_22_shiftAmt_T_2 = ans_22_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_22_shiftAmt = ans_22_expRaw > 6'h3 ? _ans_22_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_22_mantissaRaw_T = ans_22_absClipped >> ans_22_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_22_mantissaRaw = _ans_22_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_22_mantissa = ans_22_expRaw >= 6'h3 ? ans_22_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_22_expAdjusted = ans_22_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_22_exp_T_4 = ans_22_expAdjusted > 7'hf ? 4'hf : ans_22_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_22_exp = ans_22_isZero ? 4'h0 : _ans_22_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_22_fp8 = {ans_22_clippedX[31],ans_22_exp,ans_22_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_23 = {24'h0,linear_bias_23}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_23 = tempSum_23 + biasExtended_23; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_23_sign = sum32_23[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_23_absX_T = ~sum32_23; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_23_absX_T_2 = _ans_23_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_23_absX = ans_23_sign ? _ans_23_absX_T_2 : sum32_23; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_23_shiftedX_T_1 = _GEN_10432 - ans_23_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_23_shiftedX_T_3 = ans_23_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_23_shiftedX = ans_23_sign ? _ans_23_shiftedX_T_1 : _ans_23_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_23_scaledX_T_1 = ans_23_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_23_scaledX = _ans_23_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_23_clippedX_T_2 = ans_23_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_23_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_23_clippedX = ans_23_scaledX > 49'h1c0 ? 49'h1c0 : _ans_23_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_23_absClipped_T_1 = ~ans_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_23_absClipped_T_3 = _ans_23_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_23_absClipped = ans_23_clippedX[31] ? _ans_23_absClipped_T_3 : ans_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_23_isZero = ans_23_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10687 = {{16'd0}, ans_23_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_4 = _GEN_10687 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_6 = {ans_23_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_8 = _ans_23_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_9 = _ans_23_leadingZeros_T_4 | _ans_23_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10688 = {{8'd0}, _ans_23_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_14 = _GEN_10688 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_16 = {_ans_23_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_18 = _ans_23_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_19 = _ans_23_leadingZeros_T_14 | _ans_23_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10689 = {{4'd0}, _ans_23_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_24 = _GEN_10689 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_26 = {_ans_23_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_28 = _ans_23_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_29 = _ans_23_leadingZeros_T_24 | _ans_23_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10690 = {{2'd0}, _ans_23_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_34 = _GEN_10690 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_36 = {_ans_23_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_38 = _ans_23_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_39 = _ans_23_leadingZeros_T_34 | _ans_23_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10691 = {{1'd0}, _ans_23_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_44 = _GEN_10691 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_46 = {_ans_23_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_48 = _ans_23_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_23_leadingZeros_T_49 = _ans_23_leadingZeros_T_44 | _ans_23_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10692 = {{8'd0}, ans_23_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_55 = _GEN_10692 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_57 = {ans_23_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_59 = _ans_23_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_60 = _ans_23_leadingZeros_T_55 | _ans_23_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10693 = {{4'd0}, _ans_23_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_65 = _GEN_10693 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_67 = {_ans_23_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_69 = _ans_23_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_70 = _ans_23_leadingZeros_T_65 | _ans_23_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10694 = {{2'd0}, _ans_23_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_75 = _GEN_10694 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_77 = {_ans_23_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_79 = _ans_23_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_80 = _ans_23_leadingZeros_T_75 | _ans_23_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10695 = {{1'd0}, _ans_23_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_85 = _GEN_10695 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_87 = {_ans_23_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_89 = _ans_23_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_23_leadingZeros_T_90 = _ans_23_leadingZeros_T_85 | _ans_23_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_23_leadingZeros_T_93 = {_ans_23_leadingZeros_T_49,_ans_23_leadingZeros_T_90,ans_23_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_23_leadingZeros_T_143 = _ans_23_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_144 = _ans_23_leadingZeros_T_93[46] ? 6'h2e : _ans_23_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_145 = _ans_23_leadingZeros_T_93[45] ? 6'h2d : _ans_23_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_146 = _ans_23_leadingZeros_T_93[44] ? 6'h2c : _ans_23_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_147 = _ans_23_leadingZeros_T_93[43] ? 6'h2b : _ans_23_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_148 = _ans_23_leadingZeros_T_93[42] ? 6'h2a : _ans_23_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_149 = _ans_23_leadingZeros_T_93[41] ? 6'h29 : _ans_23_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_150 = _ans_23_leadingZeros_T_93[40] ? 6'h28 : _ans_23_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_151 = _ans_23_leadingZeros_T_93[39] ? 6'h27 : _ans_23_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_152 = _ans_23_leadingZeros_T_93[38] ? 6'h26 : _ans_23_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_153 = _ans_23_leadingZeros_T_93[37] ? 6'h25 : _ans_23_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_154 = _ans_23_leadingZeros_T_93[36] ? 6'h24 : _ans_23_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_155 = _ans_23_leadingZeros_T_93[35] ? 6'h23 : _ans_23_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_156 = _ans_23_leadingZeros_T_93[34] ? 6'h22 : _ans_23_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_157 = _ans_23_leadingZeros_T_93[33] ? 6'h21 : _ans_23_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_158 = _ans_23_leadingZeros_T_93[32] ? 6'h20 : _ans_23_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_159 = _ans_23_leadingZeros_T_93[31] ? 6'h1f : _ans_23_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_160 = _ans_23_leadingZeros_T_93[30] ? 6'h1e : _ans_23_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_161 = _ans_23_leadingZeros_T_93[29] ? 6'h1d : _ans_23_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_162 = _ans_23_leadingZeros_T_93[28] ? 6'h1c : _ans_23_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_163 = _ans_23_leadingZeros_T_93[27] ? 6'h1b : _ans_23_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_164 = _ans_23_leadingZeros_T_93[26] ? 6'h1a : _ans_23_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_165 = _ans_23_leadingZeros_T_93[25] ? 6'h19 : _ans_23_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_166 = _ans_23_leadingZeros_T_93[24] ? 6'h18 : _ans_23_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_167 = _ans_23_leadingZeros_T_93[23] ? 6'h17 : _ans_23_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_168 = _ans_23_leadingZeros_T_93[22] ? 6'h16 : _ans_23_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_169 = _ans_23_leadingZeros_T_93[21] ? 6'h15 : _ans_23_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_170 = _ans_23_leadingZeros_T_93[20] ? 6'h14 : _ans_23_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_171 = _ans_23_leadingZeros_T_93[19] ? 6'h13 : _ans_23_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_172 = _ans_23_leadingZeros_T_93[18] ? 6'h12 : _ans_23_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_173 = _ans_23_leadingZeros_T_93[17] ? 6'h11 : _ans_23_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_174 = _ans_23_leadingZeros_T_93[16] ? 6'h10 : _ans_23_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_175 = _ans_23_leadingZeros_T_93[15] ? 6'hf : _ans_23_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_176 = _ans_23_leadingZeros_T_93[14] ? 6'he : _ans_23_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_177 = _ans_23_leadingZeros_T_93[13] ? 6'hd : _ans_23_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_178 = _ans_23_leadingZeros_T_93[12] ? 6'hc : _ans_23_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_179 = _ans_23_leadingZeros_T_93[11] ? 6'hb : _ans_23_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_180 = _ans_23_leadingZeros_T_93[10] ? 6'ha : _ans_23_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_181 = _ans_23_leadingZeros_T_93[9] ? 6'h9 : _ans_23_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_182 = _ans_23_leadingZeros_T_93[8] ? 6'h8 : _ans_23_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_183 = _ans_23_leadingZeros_T_93[7] ? 6'h7 : _ans_23_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_184 = _ans_23_leadingZeros_T_93[6] ? 6'h6 : _ans_23_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_185 = _ans_23_leadingZeros_T_93[5] ? 6'h5 : _ans_23_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_186 = _ans_23_leadingZeros_T_93[4] ? 6'h4 : _ans_23_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_187 = _ans_23_leadingZeros_T_93[3] ? 6'h3 : _ans_23_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_188 = _ans_23_leadingZeros_T_93[2] ? 6'h2 : _ans_23_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_189 = _ans_23_leadingZeros_T_93[1] ? 6'h1 : _ans_23_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_23_leadingZeros = _ans_23_leadingZeros_T_93[0] ? 6'h0 : _ans_23_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_expRaw_T_1 = 6'h1f - ans_23_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_23_expRaw = ans_23_isZero ? 6'h0 : _ans_23_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_23_shiftAmt_T_2 = ans_23_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_23_shiftAmt = ans_23_expRaw > 6'h3 ? _ans_23_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_23_mantissaRaw_T = ans_23_absClipped >> ans_23_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_23_mantissaRaw = _ans_23_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_23_mantissa = ans_23_expRaw >= 6'h3 ? ans_23_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_23_expAdjusted = ans_23_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_23_exp_T_4 = ans_23_expAdjusted > 7'hf ? 4'hf : ans_23_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_23_exp = ans_23_isZero ? 4'h0 : _ans_23_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_23_fp8 = {ans_23_clippedX[31],ans_23_exp,ans_23_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_24 = {24'h0,linear_bias_24}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_24 = tempSum_24 + biasExtended_24; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_24_sign = sum32_24[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_24_absX_T = ~sum32_24; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_24_absX_T_2 = _ans_24_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_24_absX = ans_24_sign ? _ans_24_absX_T_2 : sum32_24; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_24_shiftedX_T_1 = _GEN_10432 - ans_24_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_24_shiftedX_T_3 = ans_24_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_24_shiftedX = ans_24_sign ? _ans_24_shiftedX_T_1 : _ans_24_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_24_scaledX_T_1 = ans_24_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_24_scaledX = _ans_24_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_24_clippedX_T_2 = ans_24_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_24_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_24_clippedX = ans_24_scaledX > 49'h1c0 ? 49'h1c0 : _ans_24_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_24_absClipped_T_1 = ~ans_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_24_absClipped_T_3 = _ans_24_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_24_absClipped = ans_24_clippedX[31] ? _ans_24_absClipped_T_3 : ans_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_24_isZero = ans_24_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10698 = {{16'd0}, ans_24_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_4 = _GEN_10698 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_6 = {ans_24_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_8 = _ans_24_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_9 = _ans_24_leadingZeros_T_4 | _ans_24_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10699 = {{8'd0}, _ans_24_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_14 = _GEN_10699 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_16 = {_ans_24_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_18 = _ans_24_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_19 = _ans_24_leadingZeros_T_14 | _ans_24_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10700 = {{4'd0}, _ans_24_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_24 = _GEN_10700 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_26 = {_ans_24_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_28 = _ans_24_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_29 = _ans_24_leadingZeros_T_24 | _ans_24_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10701 = {{2'd0}, _ans_24_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_34 = _GEN_10701 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_36 = {_ans_24_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_38 = _ans_24_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_39 = _ans_24_leadingZeros_T_34 | _ans_24_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10702 = {{1'd0}, _ans_24_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_44 = _GEN_10702 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_46 = {_ans_24_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_48 = _ans_24_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_24_leadingZeros_T_49 = _ans_24_leadingZeros_T_44 | _ans_24_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10703 = {{8'd0}, ans_24_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_55 = _GEN_10703 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_57 = {ans_24_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_59 = _ans_24_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_60 = _ans_24_leadingZeros_T_55 | _ans_24_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10704 = {{4'd0}, _ans_24_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_65 = _GEN_10704 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_67 = {_ans_24_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_69 = _ans_24_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_70 = _ans_24_leadingZeros_T_65 | _ans_24_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10705 = {{2'd0}, _ans_24_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_75 = _GEN_10705 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_77 = {_ans_24_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_79 = _ans_24_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_80 = _ans_24_leadingZeros_T_75 | _ans_24_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10706 = {{1'd0}, _ans_24_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_85 = _GEN_10706 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_87 = {_ans_24_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_89 = _ans_24_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_24_leadingZeros_T_90 = _ans_24_leadingZeros_T_85 | _ans_24_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_24_leadingZeros_T_93 = {_ans_24_leadingZeros_T_49,_ans_24_leadingZeros_T_90,ans_24_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_24_leadingZeros_T_143 = _ans_24_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_144 = _ans_24_leadingZeros_T_93[46] ? 6'h2e : _ans_24_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_145 = _ans_24_leadingZeros_T_93[45] ? 6'h2d : _ans_24_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_146 = _ans_24_leadingZeros_T_93[44] ? 6'h2c : _ans_24_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_147 = _ans_24_leadingZeros_T_93[43] ? 6'h2b : _ans_24_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_148 = _ans_24_leadingZeros_T_93[42] ? 6'h2a : _ans_24_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_149 = _ans_24_leadingZeros_T_93[41] ? 6'h29 : _ans_24_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_150 = _ans_24_leadingZeros_T_93[40] ? 6'h28 : _ans_24_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_151 = _ans_24_leadingZeros_T_93[39] ? 6'h27 : _ans_24_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_152 = _ans_24_leadingZeros_T_93[38] ? 6'h26 : _ans_24_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_153 = _ans_24_leadingZeros_T_93[37] ? 6'h25 : _ans_24_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_154 = _ans_24_leadingZeros_T_93[36] ? 6'h24 : _ans_24_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_155 = _ans_24_leadingZeros_T_93[35] ? 6'h23 : _ans_24_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_156 = _ans_24_leadingZeros_T_93[34] ? 6'h22 : _ans_24_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_157 = _ans_24_leadingZeros_T_93[33] ? 6'h21 : _ans_24_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_158 = _ans_24_leadingZeros_T_93[32] ? 6'h20 : _ans_24_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_159 = _ans_24_leadingZeros_T_93[31] ? 6'h1f : _ans_24_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_160 = _ans_24_leadingZeros_T_93[30] ? 6'h1e : _ans_24_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_161 = _ans_24_leadingZeros_T_93[29] ? 6'h1d : _ans_24_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_162 = _ans_24_leadingZeros_T_93[28] ? 6'h1c : _ans_24_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_163 = _ans_24_leadingZeros_T_93[27] ? 6'h1b : _ans_24_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_164 = _ans_24_leadingZeros_T_93[26] ? 6'h1a : _ans_24_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_165 = _ans_24_leadingZeros_T_93[25] ? 6'h19 : _ans_24_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_166 = _ans_24_leadingZeros_T_93[24] ? 6'h18 : _ans_24_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_167 = _ans_24_leadingZeros_T_93[23] ? 6'h17 : _ans_24_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_168 = _ans_24_leadingZeros_T_93[22] ? 6'h16 : _ans_24_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_169 = _ans_24_leadingZeros_T_93[21] ? 6'h15 : _ans_24_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_170 = _ans_24_leadingZeros_T_93[20] ? 6'h14 : _ans_24_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_171 = _ans_24_leadingZeros_T_93[19] ? 6'h13 : _ans_24_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_172 = _ans_24_leadingZeros_T_93[18] ? 6'h12 : _ans_24_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_173 = _ans_24_leadingZeros_T_93[17] ? 6'h11 : _ans_24_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_174 = _ans_24_leadingZeros_T_93[16] ? 6'h10 : _ans_24_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_175 = _ans_24_leadingZeros_T_93[15] ? 6'hf : _ans_24_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_176 = _ans_24_leadingZeros_T_93[14] ? 6'he : _ans_24_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_177 = _ans_24_leadingZeros_T_93[13] ? 6'hd : _ans_24_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_178 = _ans_24_leadingZeros_T_93[12] ? 6'hc : _ans_24_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_179 = _ans_24_leadingZeros_T_93[11] ? 6'hb : _ans_24_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_180 = _ans_24_leadingZeros_T_93[10] ? 6'ha : _ans_24_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_181 = _ans_24_leadingZeros_T_93[9] ? 6'h9 : _ans_24_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_182 = _ans_24_leadingZeros_T_93[8] ? 6'h8 : _ans_24_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_183 = _ans_24_leadingZeros_T_93[7] ? 6'h7 : _ans_24_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_184 = _ans_24_leadingZeros_T_93[6] ? 6'h6 : _ans_24_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_185 = _ans_24_leadingZeros_T_93[5] ? 6'h5 : _ans_24_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_186 = _ans_24_leadingZeros_T_93[4] ? 6'h4 : _ans_24_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_187 = _ans_24_leadingZeros_T_93[3] ? 6'h3 : _ans_24_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_188 = _ans_24_leadingZeros_T_93[2] ? 6'h2 : _ans_24_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_189 = _ans_24_leadingZeros_T_93[1] ? 6'h1 : _ans_24_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_24_leadingZeros = _ans_24_leadingZeros_T_93[0] ? 6'h0 : _ans_24_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_expRaw_T_1 = 6'h1f - ans_24_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_24_expRaw = ans_24_isZero ? 6'h0 : _ans_24_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_24_shiftAmt_T_2 = ans_24_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_24_shiftAmt = ans_24_expRaw > 6'h3 ? _ans_24_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_24_mantissaRaw_T = ans_24_absClipped >> ans_24_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_24_mantissaRaw = _ans_24_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_24_mantissa = ans_24_expRaw >= 6'h3 ? ans_24_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_24_expAdjusted = ans_24_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_24_exp_T_4 = ans_24_expAdjusted > 7'hf ? 4'hf : ans_24_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_24_exp = ans_24_isZero ? 4'h0 : _ans_24_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_24_fp8 = {ans_24_clippedX[31],ans_24_exp,ans_24_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_25 = {24'h0,linear_bias_25}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_25 = tempSum_25 + biasExtended_25; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_25_sign = sum32_25[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_25_absX_T = ~sum32_25; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_25_absX_T_2 = _ans_25_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_25_absX = ans_25_sign ? _ans_25_absX_T_2 : sum32_25; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_25_shiftedX_T_1 = _GEN_10432 - ans_25_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_25_shiftedX_T_3 = ans_25_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_25_shiftedX = ans_25_sign ? _ans_25_shiftedX_T_1 : _ans_25_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_25_scaledX_T_1 = ans_25_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_25_scaledX = _ans_25_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_25_clippedX_T_2 = ans_25_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_25_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_25_clippedX = ans_25_scaledX > 49'h1c0 ? 49'h1c0 : _ans_25_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_25_absClipped_T_1 = ~ans_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_25_absClipped_T_3 = _ans_25_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_25_absClipped = ans_25_clippedX[31] ? _ans_25_absClipped_T_3 : ans_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_25_isZero = ans_25_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10709 = {{16'd0}, ans_25_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_4 = _GEN_10709 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_6 = {ans_25_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_8 = _ans_25_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_9 = _ans_25_leadingZeros_T_4 | _ans_25_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10710 = {{8'd0}, _ans_25_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_14 = _GEN_10710 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_16 = {_ans_25_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_18 = _ans_25_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_19 = _ans_25_leadingZeros_T_14 | _ans_25_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10711 = {{4'd0}, _ans_25_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_24 = _GEN_10711 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_26 = {_ans_25_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_28 = _ans_25_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_29 = _ans_25_leadingZeros_T_24 | _ans_25_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10712 = {{2'd0}, _ans_25_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_34 = _GEN_10712 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_36 = {_ans_25_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_38 = _ans_25_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_39 = _ans_25_leadingZeros_T_34 | _ans_25_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10713 = {{1'd0}, _ans_25_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_44 = _GEN_10713 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_46 = {_ans_25_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_48 = _ans_25_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_25_leadingZeros_T_49 = _ans_25_leadingZeros_T_44 | _ans_25_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10714 = {{8'd0}, ans_25_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_55 = _GEN_10714 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_57 = {ans_25_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_59 = _ans_25_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_60 = _ans_25_leadingZeros_T_55 | _ans_25_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10715 = {{4'd0}, _ans_25_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_65 = _GEN_10715 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_67 = {_ans_25_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_69 = _ans_25_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_70 = _ans_25_leadingZeros_T_65 | _ans_25_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10716 = {{2'd0}, _ans_25_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_75 = _GEN_10716 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_77 = {_ans_25_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_79 = _ans_25_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_80 = _ans_25_leadingZeros_T_75 | _ans_25_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10717 = {{1'd0}, _ans_25_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_85 = _GEN_10717 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_87 = {_ans_25_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_89 = _ans_25_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_25_leadingZeros_T_90 = _ans_25_leadingZeros_T_85 | _ans_25_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_25_leadingZeros_T_93 = {_ans_25_leadingZeros_T_49,_ans_25_leadingZeros_T_90,ans_25_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_25_leadingZeros_T_143 = _ans_25_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_144 = _ans_25_leadingZeros_T_93[46] ? 6'h2e : _ans_25_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_145 = _ans_25_leadingZeros_T_93[45] ? 6'h2d : _ans_25_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_146 = _ans_25_leadingZeros_T_93[44] ? 6'h2c : _ans_25_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_147 = _ans_25_leadingZeros_T_93[43] ? 6'h2b : _ans_25_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_148 = _ans_25_leadingZeros_T_93[42] ? 6'h2a : _ans_25_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_149 = _ans_25_leadingZeros_T_93[41] ? 6'h29 : _ans_25_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_150 = _ans_25_leadingZeros_T_93[40] ? 6'h28 : _ans_25_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_151 = _ans_25_leadingZeros_T_93[39] ? 6'h27 : _ans_25_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_152 = _ans_25_leadingZeros_T_93[38] ? 6'h26 : _ans_25_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_153 = _ans_25_leadingZeros_T_93[37] ? 6'h25 : _ans_25_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_154 = _ans_25_leadingZeros_T_93[36] ? 6'h24 : _ans_25_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_155 = _ans_25_leadingZeros_T_93[35] ? 6'h23 : _ans_25_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_156 = _ans_25_leadingZeros_T_93[34] ? 6'h22 : _ans_25_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_157 = _ans_25_leadingZeros_T_93[33] ? 6'h21 : _ans_25_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_158 = _ans_25_leadingZeros_T_93[32] ? 6'h20 : _ans_25_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_159 = _ans_25_leadingZeros_T_93[31] ? 6'h1f : _ans_25_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_160 = _ans_25_leadingZeros_T_93[30] ? 6'h1e : _ans_25_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_161 = _ans_25_leadingZeros_T_93[29] ? 6'h1d : _ans_25_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_162 = _ans_25_leadingZeros_T_93[28] ? 6'h1c : _ans_25_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_163 = _ans_25_leadingZeros_T_93[27] ? 6'h1b : _ans_25_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_164 = _ans_25_leadingZeros_T_93[26] ? 6'h1a : _ans_25_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_165 = _ans_25_leadingZeros_T_93[25] ? 6'h19 : _ans_25_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_166 = _ans_25_leadingZeros_T_93[24] ? 6'h18 : _ans_25_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_167 = _ans_25_leadingZeros_T_93[23] ? 6'h17 : _ans_25_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_168 = _ans_25_leadingZeros_T_93[22] ? 6'h16 : _ans_25_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_169 = _ans_25_leadingZeros_T_93[21] ? 6'h15 : _ans_25_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_170 = _ans_25_leadingZeros_T_93[20] ? 6'h14 : _ans_25_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_171 = _ans_25_leadingZeros_T_93[19] ? 6'h13 : _ans_25_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_172 = _ans_25_leadingZeros_T_93[18] ? 6'h12 : _ans_25_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_173 = _ans_25_leadingZeros_T_93[17] ? 6'h11 : _ans_25_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_174 = _ans_25_leadingZeros_T_93[16] ? 6'h10 : _ans_25_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_175 = _ans_25_leadingZeros_T_93[15] ? 6'hf : _ans_25_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_176 = _ans_25_leadingZeros_T_93[14] ? 6'he : _ans_25_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_177 = _ans_25_leadingZeros_T_93[13] ? 6'hd : _ans_25_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_178 = _ans_25_leadingZeros_T_93[12] ? 6'hc : _ans_25_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_179 = _ans_25_leadingZeros_T_93[11] ? 6'hb : _ans_25_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_180 = _ans_25_leadingZeros_T_93[10] ? 6'ha : _ans_25_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_181 = _ans_25_leadingZeros_T_93[9] ? 6'h9 : _ans_25_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_182 = _ans_25_leadingZeros_T_93[8] ? 6'h8 : _ans_25_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_183 = _ans_25_leadingZeros_T_93[7] ? 6'h7 : _ans_25_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_184 = _ans_25_leadingZeros_T_93[6] ? 6'h6 : _ans_25_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_185 = _ans_25_leadingZeros_T_93[5] ? 6'h5 : _ans_25_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_186 = _ans_25_leadingZeros_T_93[4] ? 6'h4 : _ans_25_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_187 = _ans_25_leadingZeros_T_93[3] ? 6'h3 : _ans_25_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_188 = _ans_25_leadingZeros_T_93[2] ? 6'h2 : _ans_25_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_189 = _ans_25_leadingZeros_T_93[1] ? 6'h1 : _ans_25_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_25_leadingZeros = _ans_25_leadingZeros_T_93[0] ? 6'h0 : _ans_25_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_expRaw_T_1 = 6'h1f - ans_25_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_25_expRaw = ans_25_isZero ? 6'h0 : _ans_25_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_25_shiftAmt_T_2 = ans_25_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_25_shiftAmt = ans_25_expRaw > 6'h3 ? _ans_25_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_25_mantissaRaw_T = ans_25_absClipped >> ans_25_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_25_mantissaRaw = _ans_25_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_25_mantissa = ans_25_expRaw >= 6'h3 ? ans_25_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_25_expAdjusted = ans_25_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_25_exp_T_4 = ans_25_expAdjusted > 7'hf ? 4'hf : ans_25_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_25_exp = ans_25_isZero ? 4'h0 : _ans_25_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_25_fp8 = {ans_25_clippedX[31],ans_25_exp,ans_25_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_26 = {24'h0,linear_bias_26}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_26 = tempSum_26 + biasExtended_26; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_26_sign = sum32_26[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_26_absX_T = ~sum32_26; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_26_absX_T_2 = _ans_26_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_26_absX = ans_26_sign ? _ans_26_absX_T_2 : sum32_26; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_26_shiftedX_T_1 = _GEN_10432 - ans_26_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_26_shiftedX_T_3 = ans_26_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_26_shiftedX = ans_26_sign ? _ans_26_shiftedX_T_1 : _ans_26_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_26_scaledX_T_1 = ans_26_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_26_scaledX = _ans_26_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_26_clippedX_T_2 = ans_26_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_26_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_26_clippedX = ans_26_scaledX > 49'h1c0 ? 49'h1c0 : _ans_26_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_26_absClipped_T_1 = ~ans_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_26_absClipped_T_3 = _ans_26_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_26_absClipped = ans_26_clippedX[31] ? _ans_26_absClipped_T_3 : ans_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_26_isZero = ans_26_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10720 = {{16'd0}, ans_26_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_4 = _GEN_10720 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_6 = {ans_26_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_8 = _ans_26_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_9 = _ans_26_leadingZeros_T_4 | _ans_26_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10721 = {{8'd0}, _ans_26_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_14 = _GEN_10721 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_16 = {_ans_26_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_18 = _ans_26_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_19 = _ans_26_leadingZeros_T_14 | _ans_26_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10722 = {{4'd0}, _ans_26_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_24 = _GEN_10722 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_26 = {_ans_26_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_28 = _ans_26_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_29 = _ans_26_leadingZeros_T_24 | _ans_26_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10723 = {{2'd0}, _ans_26_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_34 = _GEN_10723 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_36 = {_ans_26_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_38 = _ans_26_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_39 = _ans_26_leadingZeros_T_34 | _ans_26_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10724 = {{1'd0}, _ans_26_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_44 = _GEN_10724 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_46 = {_ans_26_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_48 = _ans_26_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_26_leadingZeros_T_49 = _ans_26_leadingZeros_T_44 | _ans_26_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10725 = {{8'd0}, ans_26_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_55 = _GEN_10725 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_57 = {ans_26_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_59 = _ans_26_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_60 = _ans_26_leadingZeros_T_55 | _ans_26_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10726 = {{4'd0}, _ans_26_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_65 = _GEN_10726 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_67 = {_ans_26_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_69 = _ans_26_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_70 = _ans_26_leadingZeros_T_65 | _ans_26_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10727 = {{2'd0}, _ans_26_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_75 = _GEN_10727 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_77 = {_ans_26_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_79 = _ans_26_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_80 = _ans_26_leadingZeros_T_75 | _ans_26_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10728 = {{1'd0}, _ans_26_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_85 = _GEN_10728 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_87 = {_ans_26_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_89 = _ans_26_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_26_leadingZeros_T_90 = _ans_26_leadingZeros_T_85 | _ans_26_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_26_leadingZeros_T_93 = {_ans_26_leadingZeros_T_49,_ans_26_leadingZeros_T_90,ans_26_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_26_leadingZeros_T_143 = _ans_26_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_144 = _ans_26_leadingZeros_T_93[46] ? 6'h2e : _ans_26_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_145 = _ans_26_leadingZeros_T_93[45] ? 6'h2d : _ans_26_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_146 = _ans_26_leadingZeros_T_93[44] ? 6'h2c : _ans_26_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_147 = _ans_26_leadingZeros_T_93[43] ? 6'h2b : _ans_26_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_148 = _ans_26_leadingZeros_T_93[42] ? 6'h2a : _ans_26_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_149 = _ans_26_leadingZeros_T_93[41] ? 6'h29 : _ans_26_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_150 = _ans_26_leadingZeros_T_93[40] ? 6'h28 : _ans_26_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_151 = _ans_26_leadingZeros_T_93[39] ? 6'h27 : _ans_26_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_152 = _ans_26_leadingZeros_T_93[38] ? 6'h26 : _ans_26_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_153 = _ans_26_leadingZeros_T_93[37] ? 6'h25 : _ans_26_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_154 = _ans_26_leadingZeros_T_93[36] ? 6'h24 : _ans_26_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_155 = _ans_26_leadingZeros_T_93[35] ? 6'h23 : _ans_26_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_156 = _ans_26_leadingZeros_T_93[34] ? 6'h22 : _ans_26_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_157 = _ans_26_leadingZeros_T_93[33] ? 6'h21 : _ans_26_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_158 = _ans_26_leadingZeros_T_93[32] ? 6'h20 : _ans_26_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_159 = _ans_26_leadingZeros_T_93[31] ? 6'h1f : _ans_26_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_160 = _ans_26_leadingZeros_T_93[30] ? 6'h1e : _ans_26_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_161 = _ans_26_leadingZeros_T_93[29] ? 6'h1d : _ans_26_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_162 = _ans_26_leadingZeros_T_93[28] ? 6'h1c : _ans_26_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_163 = _ans_26_leadingZeros_T_93[27] ? 6'h1b : _ans_26_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_164 = _ans_26_leadingZeros_T_93[26] ? 6'h1a : _ans_26_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_165 = _ans_26_leadingZeros_T_93[25] ? 6'h19 : _ans_26_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_166 = _ans_26_leadingZeros_T_93[24] ? 6'h18 : _ans_26_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_167 = _ans_26_leadingZeros_T_93[23] ? 6'h17 : _ans_26_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_168 = _ans_26_leadingZeros_T_93[22] ? 6'h16 : _ans_26_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_169 = _ans_26_leadingZeros_T_93[21] ? 6'h15 : _ans_26_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_170 = _ans_26_leadingZeros_T_93[20] ? 6'h14 : _ans_26_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_171 = _ans_26_leadingZeros_T_93[19] ? 6'h13 : _ans_26_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_172 = _ans_26_leadingZeros_T_93[18] ? 6'h12 : _ans_26_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_173 = _ans_26_leadingZeros_T_93[17] ? 6'h11 : _ans_26_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_174 = _ans_26_leadingZeros_T_93[16] ? 6'h10 : _ans_26_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_175 = _ans_26_leadingZeros_T_93[15] ? 6'hf : _ans_26_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_176 = _ans_26_leadingZeros_T_93[14] ? 6'he : _ans_26_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_177 = _ans_26_leadingZeros_T_93[13] ? 6'hd : _ans_26_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_178 = _ans_26_leadingZeros_T_93[12] ? 6'hc : _ans_26_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_179 = _ans_26_leadingZeros_T_93[11] ? 6'hb : _ans_26_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_180 = _ans_26_leadingZeros_T_93[10] ? 6'ha : _ans_26_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_181 = _ans_26_leadingZeros_T_93[9] ? 6'h9 : _ans_26_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_182 = _ans_26_leadingZeros_T_93[8] ? 6'h8 : _ans_26_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_183 = _ans_26_leadingZeros_T_93[7] ? 6'h7 : _ans_26_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_184 = _ans_26_leadingZeros_T_93[6] ? 6'h6 : _ans_26_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_185 = _ans_26_leadingZeros_T_93[5] ? 6'h5 : _ans_26_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_186 = _ans_26_leadingZeros_T_93[4] ? 6'h4 : _ans_26_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_187 = _ans_26_leadingZeros_T_93[3] ? 6'h3 : _ans_26_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_188 = _ans_26_leadingZeros_T_93[2] ? 6'h2 : _ans_26_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_189 = _ans_26_leadingZeros_T_93[1] ? 6'h1 : _ans_26_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_26_leadingZeros = _ans_26_leadingZeros_T_93[0] ? 6'h0 : _ans_26_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_expRaw_T_1 = 6'h1f - ans_26_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_26_expRaw = ans_26_isZero ? 6'h0 : _ans_26_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_26_shiftAmt_T_2 = ans_26_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_26_shiftAmt = ans_26_expRaw > 6'h3 ? _ans_26_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_26_mantissaRaw_T = ans_26_absClipped >> ans_26_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_26_mantissaRaw = _ans_26_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_26_mantissa = ans_26_expRaw >= 6'h3 ? ans_26_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_26_expAdjusted = ans_26_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_26_exp_T_4 = ans_26_expAdjusted > 7'hf ? 4'hf : ans_26_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_26_exp = ans_26_isZero ? 4'h0 : _ans_26_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_26_fp8 = {ans_26_clippedX[31],ans_26_exp,ans_26_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_27 = {24'h0,linear_bias_27}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_27 = tempSum_27 + biasExtended_27; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_27_sign = sum32_27[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_27_absX_T = ~sum32_27; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_27_absX_T_2 = _ans_27_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_27_absX = ans_27_sign ? _ans_27_absX_T_2 : sum32_27; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_27_shiftedX_T_1 = _GEN_10432 - ans_27_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_27_shiftedX_T_3 = ans_27_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_27_shiftedX = ans_27_sign ? _ans_27_shiftedX_T_1 : _ans_27_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_27_scaledX_T_1 = ans_27_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_27_scaledX = _ans_27_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_27_clippedX_T_2 = ans_27_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_27_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_27_clippedX = ans_27_scaledX > 49'h1c0 ? 49'h1c0 : _ans_27_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_27_absClipped_T_1 = ~ans_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_27_absClipped_T_3 = _ans_27_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_27_absClipped = ans_27_clippedX[31] ? _ans_27_absClipped_T_3 : ans_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_27_isZero = ans_27_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10731 = {{16'd0}, ans_27_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_4 = _GEN_10731 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_6 = {ans_27_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_8 = _ans_27_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_9 = _ans_27_leadingZeros_T_4 | _ans_27_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10732 = {{8'd0}, _ans_27_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_14 = _GEN_10732 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_16 = {_ans_27_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_18 = _ans_27_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_19 = _ans_27_leadingZeros_T_14 | _ans_27_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10733 = {{4'd0}, _ans_27_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_24 = _GEN_10733 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_26 = {_ans_27_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_28 = _ans_27_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_29 = _ans_27_leadingZeros_T_24 | _ans_27_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10734 = {{2'd0}, _ans_27_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_34 = _GEN_10734 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_36 = {_ans_27_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_38 = _ans_27_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_39 = _ans_27_leadingZeros_T_34 | _ans_27_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10735 = {{1'd0}, _ans_27_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_44 = _GEN_10735 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_46 = {_ans_27_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_48 = _ans_27_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_27_leadingZeros_T_49 = _ans_27_leadingZeros_T_44 | _ans_27_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10736 = {{8'd0}, ans_27_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_55 = _GEN_10736 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_57 = {ans_27_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_59 = _ans_27_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_60 = _ans_27_leadingZeros_T_55 | _ans_27_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10737 = {{4'd0}, _ans_27_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_65 = _GEN_10737 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_67 = {_ans_27_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_69 = _ans_27_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_70 = _ans_27_leadingZeros_T_65 | _ans_27_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10738 = {{2'd0}, _ans_27_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_75 = _GEN_10738 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_77 = {_ans_27_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_79 = _ans_27_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_80 = _ans_27_leadingZeros_T_75 | _ans_27_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10739 = {{1'd0}, _ans_27_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_85 = _GEN_10739 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_87 = {_ans_27_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_89 = _ans_27_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_27_leadingZeros_T_90 = _ans_27_leadingZeros_T_85 | _ans_27_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_27_leadingZeros_T_93 = {_ans_27_leadingZeros_T_49,_ans_27_leadingZeros_T_90,ans_27_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_27_leadingZeros_T_143 = _ans_27_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_144 = _ans_27_leadingZeros_T_93[46] ? 6'h2e : _ans_27_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_145 = _ans_27_leadingZeros_T_93[45] ? 6'h2d : _ans_27_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_146 = _ans_27_leadingZeros_T_93[44] ? 6'h2c : _ans_27_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_147 = _ans_27_leadingZeros_T_93[43] ? 6'h2b : _ans_27_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_148 = _ans_27_leadingZeros_T_93[42] ? 6'h2a : _ans_27_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_149 = _ans_27_leadingZeros_T_93[41] ? 6'h29 : _ans_27_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_150 = _ans_27_leadingZeros_T_93[40] ? 6'h28 : _ans_27_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_151 = _ans_27_leadingZeros_T_93[39] ? 6'h27 : _ans_27_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_152 = _ans_27_leadingZeros_T_93[38] ? 6'h26 : _ans_27_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_153 = _ans_27_leadingZeros_T_93[37] ? 6'h25 : _ans_27_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_154 = _ans_27_leadingZeros_T_93[36] ? 6'h24 : _ans_27_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_155 = _ans_27_leadingZeros_T_93[35] ? 6'h23 : _ans_27_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_156 = _ans_27_leadingZeros_T_93[34] ? 6'h22 : _ans_27_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_157 = _ans_27_leadingZeros_T_93[33] ? 6'h21 : _ans_27_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_158 = _ans_27_leadingZeros_T_93[32] ? 6'h20 : _ans_27_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_159 = _ans_27_leadingZeros_T_93[31] ? 6'h1f : _ans_27_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_160 = _ans_27_leadingZeros_T_93[30] ? 6'h1e : _ans_27_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_161 = _ans_27_leadingZeros_T_93[29] ? 6'h1d : _ans_27_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_162 = _ans_27_leadingZeros_T_93[28] ? 6'h1c : _ans_27_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_163 = _ans_27_leadingZeros_T_93[27] ? 6'h1b : _ans_27_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_164 = _ans_27_leadingZeros_T_93[26] ? 6'h1a : _ans_27_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_165 = _ans_27_leadingZeros_T_93[25] ? 6'h19 : _ans_27_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_166 = _ans_27_leadingZeros_T_93[24] ? 6'h18 : _ans_27_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_167 = _ans_27_leadingZeros_T_93[23] ? 6'h17 : _ans_27_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_168 = _ans_27_leadingZeros_T_93[22] ? 6'h16 : _ans_27_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_169 = _ans_27_leadingZeros_T_93[21] ? 6'h15 : _ans_27_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_170 = _ans_27_leadingZeros_T_93[20] ? 6'h14 : _ans_27_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_171 = _ans_27_leadingZeros_T_93[19] ? 6'h13 : _ans_27_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_172 = _ans_27_leadingZeros_T_93[18] ? 6'h12 : _ans_27_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_173 = _ans_27_leadingZeros_T_93[17] ? 6'h11 : _ans_27_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_174 = _ans_27_leadingZeros_T_93[16] ? 6'h10 : _ans_27_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_175 = _ans_27_leadingZeros_T_93[15] ? 6'hf : _ans_27_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_176 = _ans_27_leadingZeros_T_93[14] ? 6'he : _ans_27_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_177 = _ans_27_leadingZeros_T_93[13] ? 6'hd : _ans_27_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_178 = _ans_27_leadingZeros_T_93[12] ? 6'hc : _ans_27_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_179 = _ans_27_leadingZeros_T_93[11] ? 6'hb : _ans_27_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_180 = _ans_27_leadingZeros_T_93[10] ? 6'ha : _ans_27_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_181 = _ans_27_leadingZeros_T_93[9] ? 6'h9 : _ans_27_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_182 = _ans_27_leadingZeros_T_93[8] ? 6'h8 : _ans_27_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_183 = _ans_27_leadingZeros_T_93[7] ? 6'h7 : _ans_27_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_184 = _ans_27_leadingZeros_T_93[6] ? 6'h6 : _ans_27_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_185 = _ans_27_leadingZeros_T_93[5] ? 6'h5 : _ans_27_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_186 = _ans_27_leadingZeros_T_93[4] ? 6'h4 : _ans_27_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_187 = _ans_27_leadingZeros_T_93[3] ? 6'h3 : _ans_27_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_188 = _ans_27_leadingZeros_T_93[2] ? 6'h2 : _ans_27_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_189 = _ans_27_leadingZeros_T_93[1] ? 6'h1 : _ans_27_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_27_leadingZeros = _ans_27_leadingZeros_T_93[0] ? 6'h0 : _ans_27_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_expRaw_T_1 = 6'h1f - ans_27_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_27_expRaw = ans_27_isZero ? 6'h0 : _ans_27_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_27_shiftAmt_T_2 = ans_27_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_27_shiftAmt = ans_27_expRaw > 6'h3 ? _ans_27_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_27_mantissaRaw_T = ans_27_absClipped >> ans_27_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_27_mantissaRaw = _ans_27_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_27_mantissa = ans_27_expRaw >= 6'h3 ? ans_27_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_27_expAdjusted = ans_27_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_27_exp_T_4 = ans_27_expAdjusted > 7'hf ? 4'hf : ans_27_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_27_exp = ans_27_isZero ? 4'h0 : _ans_27_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_27_fp8 = {ans_27_clippedX[31],ans_27_exp,ans_27_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_28 = {24'h0,linear_bias_28}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_28 = tempSum_28 + biasExtended_28; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_28_sign = sum32_28[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_28_absX_T = ~sum32_28; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_28_absX_T_2 = _ans_28_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_28_absX = ans_28_sign ? _ans_28_absX_T_2 : sum32_28; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_28_shiftedX_T_1 = _GEN_10432 - ans_28_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_28_shiftedX_T_3 = ans_28_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_28_shiftedX = ans_28_sign ? _ans_28_shiftedX_T_1 : _ans_28_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_28_scaledX_T_1 = ans_28_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_28_scaledX = _ans_28_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_28_clippedX_T_2 = ans_28_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_28_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_28_clippedX = ans_28_scaledX > 49'h1c0 ? 49'h1c0 : _ans_28_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_28_absClipped_T_1 = ~ans_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_28_absClipped_T_3 = _ans_28_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_28_absClipped = ans_28_clippedX[31] ? _ans_28_absClipped_T_3 : ans_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_28_isZero = ans_28_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10742 = {{16'd0}, ans_28_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_4 = _GEN_10742 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_6 = {ans_28_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_8 = _ans_28_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_9 = _ans_28_leadingZeros_T_4 | _ans_28_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10743 = {{8'd0}, _ans_28_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_14 = _GEN_10743 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_16 = {_ans_28_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_18 = _ans_28_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_19 = _ans_28_leadingZeros_T_14 | _ans_28_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10744 = {{4'd0}, _ans_28_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_24 = _GEN_10744 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_26 = {_ans_28_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_28 = _ans_28_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_29 = _ans_28_leadingZeros_T_24 | _ans_28_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10745 = {{2'd0}, _ans_28_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_34 = _GEN_10745 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_36 = {_ans_28_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_38 = _ans_28_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_39 = _ans_28_leadingZeros_T_34 | _ans_28_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10746 = {{1'd0}, _ans_28_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_44 = _GEN_10746 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_46 = {_ans_28_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_48 = _ans_28_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_28_leadingZeros_T_49 = _ans_28_leadingZeros_T_44 | _ans_28_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10747 = {{8'd0}, ans_28_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_55 = _GEN_10747 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_57 = {ans_28_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_59 = _ans_28_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_60 = _ans_28_leadingZeros_T_55 | _ans_28_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10748 = {{4'd0}, _ans_28_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_65 = _GEN_10748 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_67 = {_ans_28_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_69 = _ans_28_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_70 = _ans_28_leadingZeros_T_65 | _ans_28_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10749 = {{2'd0}, _ans_28_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_75 = _GEN_10749 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_77 = {_ans_28_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_79 = _ans_28_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_80 = _ans_28_leadingZeros_T_75 | _ans_28_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10750 = {{1'd0}, _ans_28_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_85 = _GEN_10750 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_87 = {_ans_28_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_89 = _ans_28_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_28_leadingZeros_T_90 = _ans_28_leadingZeros_T_85 | _ans_28_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_28_leadingZeros_T_93 = {_ans_28_leadingZeros_T_49,_ans_28_leadingZeros_T_90,ans_28_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_28_leadingZeros_T_143 = _ans_28_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_144 = _ans_28_leadingZeros_T_93[46] ? 6'h2e : _ans_28_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_145 = _ans_28_leadingZeros_T_93[45] ? 6'h2d : _ans_28_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_146 = _ans_28_leadingZeros_T_93[44] ? 6'h2c : _ans_28_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_147 = _ans_28_leadingZeros_T_93[43] ? 6'h2b : _ans_28_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_148 = _ans_28_leadingZeros_T_93[42] ? 6'h2a : _ans_28_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_149 = _ans_28_leadingZeros_T_93[41] ? 6'h29 : _ans_28_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_150 = _ans_28_leadingZeros_T_93[40] ? 6'h28 : _ans_28_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_151 = _ans_28_leadingZeros_T_93[39] ? 6'h27 : _ans_28_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_152 = _ans_28_leadingZeros_T_93[38] ? 6'h26 : _ans_28_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_153 = _ans_28_leadingZeros_T_93[37] ? 6'h25 : _ans_28_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_154 = _ans_28_leadingZeros_T_93[36] ? 6'h24 : _ans_28_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_155 = _ans_28_leadingZeros_T_93[35] ? 6'h23 : _ans_28_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_156 = _ans_28_leadingZeros_T_93[34] ? 6'h22 : _ans_28_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_157 = _ans_28_leadingZeros_T_93[33] ? 6'h21 : _ans_28_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_158 = _ans_28_leadingZeros_T_93[32] ? 6'h20 : _ans_28_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_159 = _ans_28_leadingZeros_T_93[31] ? 6'h1f : _ans_28_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_160 = _ans_28_leadingZeros_T_93[30] ? 6'h1e : _ans_28_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_161 = _ans_28_leadingZeros_T_93[29] ? 6'h1d : _ans_28_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_162 = _ans_28_leadingZeros_T_93[28] ? 6'h1c : _ans_28_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_163 = _ans_28_leadingZeros_T_93[27] ? 6'h1b : _ans_28_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_164 = _ans_28_leadingZeros_T_93[26] ? 6'h1a : _ans_28_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_165 = _ans_28_leadingZeros_T_93[25] ? 6'h19 : _ans_28_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_166 = _ans_28_leadingZeros_T_93[24] ? 6'h18 : _ans_28_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_167 = _ans_28_leadingZeros_T_93[23] ? 6'h17 : _ans_28_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_168 = _ans_28_leadingZeros_T_93[22] ? 6'h16 : _ans_28_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_169 = _ans_28_leadingZeros_T_93[21] ? 6'h15 : _ans_28_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_170 = _ans_28_leadingZeros_T_93[20] ? 6'h14 : _ans_28_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_171 = _ans_28_leadingZeros_T_93[19] ? 6'h13 : _ans_28_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_172 = _ans_28_leadingZeros_T_93[18] ? 6'h12 : _ans_28_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_173 = _ans_28_leadingZeros_T_93[17] ? 6'h11 : _ans_28_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_174 = _ans_28_leadingZeros_T_93[16] ? 6'h10 : _ans_28_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_175 = _ans_28_leadingZeros_T_93[15] ? 6'hf : _ans_28_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_176 = _ans_28_leadingZeros_T_93[14] ? 6'he : _ans_28_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_177 = _ans_28_leadingZeros_T_93[13] ? 6'hd : _ans_28_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_178 = _ans_28_leadingZeros_T_93[12] ? 6'hc : _ans_28_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_179 = _ans_28_leadingZeros_T_93[11] ? 6'hb : _ans_28_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_180 = _ans_28_leadingZeros_T_93[10] ? 6'ha : _ans_28_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_181 = _ans_28_leadingZeros_T_93[9] ? 6'h9 : _ans_28_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_182 = _ans_28_leadingZeros_T_93[8] ? 6'h8 : _ans_28_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_183 = _ans_28_leadingZeros_T_93[7] ? 6'h7 : _ans_28_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_184 = _ans_28_leadingZeros_T_93[6] ? 6'h6 : _ans_28_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_185 = _ans_28_leadingZeros_T_93[5] ? 6'h5 : _ans_28_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_186 = _ans_28_leadingZeros_T_93[4] ? 6'h4 : _ans_28_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_187 = _ans_28_leadingZeros_T_93[3] ? 6'h3 : _ans_28_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_188 = _ans_28_leadingZeros_T_93[2] ? 6'h2 : _ans_28_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_189 = _ans_28_leadingZeros_T_93[1] ? 6'h1 : _ans_28_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_28_leadingZeros = _ans_28_leadingZeros_T_93[0] ? 6'h0 : _ans_28_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_expRaw_T_1 = 6'h1f - ans_28_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_28_expRaw = ans_28_isZero ? 6'h0 : _ans_28_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_28_shiftAmt_T_2 = ans_28_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_28_shiftAmt = ans_28_expRaw > 6'h3 ? _ans_28_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_28_mantissaRaw_T = ans_28_absClipped >> ans_28_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_28_mantissaRaw = _ans_28_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_28_mantissa = ans_28_expRaw >= 6'h3 ? ans_28_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_28_expAdjusted = ans_28_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_28_exp_T_4 = ans_28_expAdjusted > 7'hf ? 4'hf : ans_28_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_28_exp = ans_28_isZero ? 4'h0 : _ans_28_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_28_fp8 = {ans_28_clippedX[31],ans_28_exp,ans_28_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_29 = {24'h0,linear_bias_29}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_29 = tempSum_29 + biasExtended_29; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_29_sign = sum32_29[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_29_absX_T = ~sum32_29; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_29_absX_T_2 = _ans_29_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_29_absX = ans_29_sign ? _ans_29_absX_T_2 : sum32_29; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_29_shiftedX_T_1 = _GEN_10432 - ans_29_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_29_shiftedX_T_3 = ans_29_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_29_shiftedX = ans_29_sign ? _ans_29_shiftedX_T_1 : _ans_29_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_29_scaledX_T_1 = ans_29_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_29_scaledX = _ans_29_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_29_clippedX_T_2 = ans_29_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_29_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_29_clippedX = ans_29_scaledX > 49'h1c0 ? 49'h1c0 : _ans_29_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_29_absClipped_T_1 = ~ans_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_29_absClipped_T_3 = _ans_29_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_29_absClipped = ans_29_clippedX[31] ? _ans_29_absClipped_T_3 : ans_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_29_isZero = ans_29_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10753 = {{16'd0}, ans_29_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_4 = _GEN_10753 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_6 = {ans_29_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_8 = _ans_29_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_9 = _ans_29_leadingZeros_T_4 | _ans_29_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10754 = {{8'd0}, _ans_29_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_14 = _GEN_10754 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_16 = {_ans_29_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_18 = _ans_29_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_19 = _ans_29_leadingZeros_T_14 | _ans_29_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10755 = {{4'd0}, _ans_29_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_24 = _GEN_10755 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_26 = {_ans_29_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_28 = _ans_29_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_29 = _ans_29_leadingZeros_T_24 | _ans_29_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10756 = {{2'd0}, _ans_29_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_34 = _GEN_10756 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_36 = {_ans_29_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_38 = _ans_29_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_39 = _ans_29_leadingZeros_T_34 | _ans_29_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10757 = {{1'd0}, _ans_29_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_44 = _GEN_10757 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_46 = {_ans_29_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_48 = _ans_29_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_29_leadingZeros_T_49 = _ans_29_leadingZeros_T_44 | _ans_29_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10758 = {{8'd0}, ans_29_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_55 = _GEN_10758 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_57 = {ans_29_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_59 = _ans_29_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_60 = _ans_29_leadingZeros_T_55 | _ans_29_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10759 = {{4'd0}, _ans_29_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_65 = _GEN_10759 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_67 = {_ans_29_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_69 = _ans_29_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_70 = _ans_29_leadingZeros_T_65 | _ans_29_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10760 = {{2'd0}, _ans_29_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_75 = _GEN_10760 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_77 = {_ans_29_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_79 = _ans_29_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_80 = _ans_29_leadingZeros_T_75 | _ans_29_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10761 = {{1'd0}, _ans_29_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_85 = _GEN_10761 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_87 = {_ans_29_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_89 = _ans_29_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_29_leadingZeros_T_90 = _ans_29_leadingZeros_T_85 | _ans_29_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_29_leadingZeros_T_93 = {_ans_29_leadingZeros_T_49,_ans_29_leadingZeros_T_90,ans_29_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_29_leadingZeros_T_143 = _ans_29_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_144 = _ans_29_leadingZeros_T_93[46] ? 6'h2e : _ans_29_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_145 = _ans_29_leadingZeros_T_93[45] ? 6'h2d : _ans_29_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_146 = _ans_29_leadingZeros_T_93[44] ? 6'h2c : _ans_29_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_147 = _ans_29_leadingZeros_T_93[43] ? 6'h2b : _ans_29_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_148 = _ans_29_leadingZeros_T_93[42] ? 6'h2a : _ans_29_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_149 = _ans_29_leadingZeros_T_93[41] ? 6'h29 : _ans_29_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_150 = _ans_29_leadingZeros_T_93[40] ? 6'h28 : _ans_29_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_151 = _ans_29_leadingZeros_T_93[39] ? 6'h27 : _ans_29_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_152 = _ans_29_leadingZeros_T_93[38] ? 6'h26 : _ans_29_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_153 = _ans_29_leadingZeros_T_93[37] ? 6'h25 : _ans_29_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_154 = _ans_29_leadingZeros_T_93[36] ? 6'h24 : _ans_29_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_155 = _ans_29_leadingZeros_T_93[35] ? 6'h23 : _ans_29_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_156 = _ans_29_leadingZeros_T_93[34] ? 6'h22 : _ans_29_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_157 = _ans_29_leadingZeros_T_93[33] ? 6'h21 : _ans_29_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_158 = _ans_29_leadingZeros_T_93[32] ? 6'h20 : _ans_29_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_159 = _ans_29_leadingZeros_T_93[31] ? 6'h1f : _ans_29_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_160 = _ans_29_leadingZeros_T_93[30] ? 6'h1e : _ans_29_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_161 = _ans_29_leadingZeros_T_93[29] ? 6'h1d : _ans_29_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_162 = _ans_29_leadingZeros_T_93[28] ? 6'h1c : _ans_29_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_163 = _ans_29_leadingZeros_T_93[27] ? 6'h1b : _ans_29_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_164 = _ans_29_leadingZeros_T_93[26] ? 6'h1a : _ans_29_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_165 = _ans_29_leadingZeros_T_93[25] ? 6'h19 : _ans_29_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_166 = _ans_29_leadingZeros_T_93[24] ? 6'h18 : _ans_29_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_167 = _ans_29_leadingZeros_T_93[23] ? 6'h17 : _ans_29_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_168 = _ans_29_leadingZeros_T_93[22] ? 6'h16 : _ans_29_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_169 = _ans_29_leadingZeros_T_93[21] ? 6'h15 : _ans_29_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_170 = _ans_29_leadingZeros_T_93[20] ? 6'h14 : _ans_29_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_171 = _ans_29_leadingZeros_T_93[19] ? 6'h13 : _ans_29_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_172 = _ans_29_leadingZeros_T_93[18] ? 6'h12 : _ans_29_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_173 = _ans_29_leadingZeros_T_93[17] ? 6'h11 : _ans_29_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_174 = _ans_29_leadingZeros_T_93[16] ? 6'h10 : _ans_29_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_175 = _ans_29_leadingZeros_T_93[15] ? 6'hf : _ans_29_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_176 = _ans_29_leadingZeros_T_93[14] ? 6'he : _ans_29_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_177 = _ans_29_leadingZeros_T_93[13] ? 6'hd : _ans_29_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_178 = _ans_29_leadingZeros_T_93[12] ? 6'hc : _ans_29_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_179 = _ans_29_leadingZeros_T_93[11] ? 6'hb : _ans_29_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_180 = _ans_29_leadingZeros_T_93[10] ? 6'ha : _ans_29_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_181 = _ans_29_leadingZeros_T_93[9] ? 6'h9 : _ans_29_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_182 = _ans_29_leadingZeros_T_93[8] ? 6'h8 : _ans_29_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_183 = _ans_29_leadingZeros_T_93[7] ? 6'h7 : _ans_29_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_184 = _ans_29_leadingZeros_T_93[6] ? 6'h6 : _ans_29_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_185 = _ans_29_leadingZeros_T_93[5] ? 6'h5 : _ans_29_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_186 = _ans_29_leadingZeros_T_93[4] ? 6'h4 : _ans_29_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_187 = _ans_29_leadingZeros_T_93[3] ? 6'h3 : _ans_29_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_188 = _ans_29_leadingZeros_T_93[2] ? 6'h2 : _ans_29_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_189 = _ans_29_leadingZeros_T_93[1] ? 6'h1 : _ans_29_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_29_leadingZeros = _ans_29_leadingZeros_T_93[0] ? 6'h0 : _ans_29_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_expRaw_T_1 = 6'h1f - ans_29_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_29_expRaw = ans_29_isZero ? 6'h0 : _ans_29_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_29_shiftAmt_T_2 = ans_29_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_29_shiftAmt = ans_29_expRaw > 6'h3 ? _ans_29_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_29_mantissaRaw_T = ans_29_absClipped >> ans_29_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_29_mantissaRaw = _ans_29_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_29_mantissa = ans_29_expRaw >= 6'h3 ? ans_29_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_29_expAdjusted = ans_29_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_29_exp_T_4 = ans_29_expAdjusted > 7'hf ? 4'hf : ans_29_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_29_exp = ans_29_isZero ? 4'h0 : _ans_29_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_29_fp8 = {ans_29_clippedX[31],ans_29_exp,ans_29_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_30 = {24'h0,linear_bias_30}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_30 = tempSum_30 + biasExtended_30; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_30_sign = sum32_30[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_30_absX_T = ~sum32_30; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_30_absX_T_2 = _ans_30_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_30_absX = ans_30_sign ? _ans_30_absX_T_2 : sum32_30; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_30_shiftedX_T_1 = _GEN_10432 - ans_30_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_30_shiftedX_T_3 = ans_30_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_30_shiftedX = ans_30_sign ? _ans_30_shiftedX_T_1 : _ans_30_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_30_scaledX_T_1 = ans_30_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_30_scaledX = _ans_30_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_30_clippedX_T_2 = ans_30_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_30_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_30_clippedX = ans_30_scaledX > 49'h1c0 ? 49'h1c0 : _ans_30_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_30_absClipped_T_1 = ~ans_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_30_absClipped_T_3 = _ans_30_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_30_absClipped = ans_30_clippedX[31] ? _ans_30_absClipped_T_3 : ans_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_30_isZero = ans_30_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10764 = {{16'd0}, ans_30_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_4 = _GEN_10764 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_6 = {ans_30_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_8 = _ans_30_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_9 = _ans_30_leadingZeros_T_4 | _ans_30_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10765 = {{8'd0}, _ans_30_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_14 = _GEN_10765 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_16 = {_ans_30_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_18 = _ans_30_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_19 = _ans_30_leadingZeros_T_14 | _ans_30_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10766 = {{4'd0}, _ans_30_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_24 = _GEN_10766 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_26 = {_ans_30_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_28 = _ans_30_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_29 = _ans_30_leadingZeros_T_24 | _ans_30_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10767 = {{2'd0}, _ans_30_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_34 = _GEN_10767 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_36 = {_ans_30_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_38 = _ans_30_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_39 = _ans_30_leadingZeros_T_34 | _ans_30_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10768 = {{1'd0}, _ans_30_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_44 = _GEN_10768 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_46 = {_ans_30_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_48 = _ans_30_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_30_leadingZeros_T_49 = _ans_30_leadingZeros_T_44 | _ans_30_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10769 = {{8'd0}, ans_30_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_55 = _GEN_10769 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_57 = {ans_30_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_59 = _ans_30_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_60 = _ans_30_leadingZeros_T_55 | _ans_30_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10770 = {{4'd0}, _ans_30_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_65 = _GEN_10770 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_67 = {_ans_30_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_69 = _ans_30_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_70 = _ans_30_leadingZeros_T_65 | _ans_30_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10771 = {{2'd0}, _ans_30_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_75 = _GEN_10771 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_77 = {_ans_30_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_79 = _ans_30_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_80 = _ans_30_leadingZeros_T_75 | _ans_30_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10772 = {{1'd0}, _ans_30_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_85 = _GEN_10772 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_87 = {_ans_30_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_89 = _ans_30_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_30_leadingZeros_T_90 = _ans_30_leadingZeros_T_85 | _ans_30_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_30_leadingZeros_T_93 = {_ans_30_leadingZeros_T_49,_ans_30_leadingZeros_T_90,ans_30_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_30_leadingZeros_T_143 = _ans_30_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_144 = _ans_30_leadingZeros_T_93[46] ? 6'h2e : _ans_30_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_145 = _ans_30_leadingZeros_T_93[45] ? 6'h2d : _ans_30_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_146 = _ans_30_leadingZeros_T_93[44] ? 6'h2c : _ans_30_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_147 = _ans_30_leadingZeros_T_93[43] ? 6'h2b : _ans_30_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_148 = _ans_30_leadingZeros_T_93[42] ? 6'h2a : _ans_30_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_149 = _ans_30_leadingZeros_T_93[41] ? 6'h29 : _ans_30_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_150 = _ans_30_leadingZeros_T_93[40] ? 6'h28 : _ans_30_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_151 = _ans_30_leadingZeros_T_93[39] ? 6'h27 : _ans_30_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_152 = _ans_30_leadingZeros_T_93[38] ? 6'h26 : _ans_30_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_153 = _ans_30_leadingZeros_T_93[37] ? 6'h25 : _ans_30_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_154 = _ans_30_leadingZeros_T_93[36] ? 6'h24 : _ans_30_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_155 = _ans_30_leadingZeros_T_93[35] ? 6'h23 : _ans_30_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_156 = _ans_30_leadingZeros_T_93[34] ? 6'h22 : _ans_30_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_157 = _ans_30_leadingZeros_T_93[33] ? 6'h21 : _ans_30_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_158 = _ans_30_leadingZeros_T_93[32] ? 6'h20 : _ans_30_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_159 = _ans_30_leadingZeros_T_93[31] ? 6'h1f : _ans_30_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_160 = _ans_30_leadingZeros_T_93[30] ? 6'h1e : _ans_30_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_161 = _ans_30_leadingZeros_T_93[29] ? 6'h1d : _ans_30_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_162 = _ans_30_leadingZeros_T_93[28] ? 6'h1c : _ans_30_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_163 = _ans_30_leadingZeros_T_93[27] ? 6'h1b : _ans_30_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_164 = _ans_30_leadingZeros_T_93[26] ? 6'h1a : _ans_30_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_165 = _ans_30_leadingZeros_T_93[25] ? 6'h19 : _ans_30_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_166 = _ans_30_leadingZeros_T_93[24] ? 6'h18 : _ans_30_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_167 = _ans_30_leadingZeros_T_93[23] ? 6'h17 : _ans_30_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_168 = _ans_30_leadingZeros_T_93[22] ? 6'h16 : _ans_30_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_169 = _ans_30_leadingZeros_T_93[21] ? 6'h15 : _ans_30_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_170 = _ans_30_leadingZeros_T_93[20] ? 6'h14 : _ans_30_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_171 = _ans_30_leadingZeros_T_93[19] ? 6'h13 : _ans_30_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_172 = _ans_30_leadingZeros_T_93[18] ? 6'h12 : _ans_30_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_173 = _ans_30_leadingZeros_T_93[17] ? 6'h11 : _ans_30_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_174 = _ans_30_leadingZeros_T_93[16] ? 6'h10 : _ans_30_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_175 = _ans_30_leadingZeros_T_93[15] ? 6'hf : _ans_30_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_176 = _ans_30_leadingZeros_T_93[14] ? 6'he : _ans_30_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_177 = _ans_30_leadingZeros_T_93[13] ? 6'hd : _ans_30_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_178 = _ans_30_leadingZeros_T_93[12] ? 6'hc : _ans_30_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_179 = _ans_30_leadingZeros_T_93[11] ? 6'hb : _ans_30_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_180 = _ans_30_leadingZeros_T_93[10] ? 6'ha : _ans_30_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_181 = _ans_30_leadingZeros_T_93[9] ? 6'h9 : _ans_30_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_182 = _ans_30_leadingZeros_T_93[8] ? 6'h8 : _ans_30_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_183 = _ans_30_leadingZeros_T_93[7] ? 6'h7 : _ans_30_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_184 = _ans_30_leadingZeros_T_93[6] ? 6'h6 : _ans_30_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_185 = _ans_30_leadingZeros_T_93[5] ? 6'h5 : _ans_30_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_186 = _ans_30_leadingZeros_T_93[4] ? 6'h4 : _ans_30_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_187 = _ans_30_leadingZeros_T_93[3] ? 6'h3 : _ans_30_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_188 = _ans_30_leadingZeros_T_93[2] ? 6'h2 : _ans_30_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_189 = _ans_30_leadingZeros_T_93[1] ? 6'h1 : _ans_30_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_30_leadingZeros = _ans_30_leadingZeros_T_93[0] ? 6'h0 : _ans_30_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_expRaw_T_1 = 6'h1f - ans_30_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_30_expRaw = ans_30_isZero ? 6'h0 : _ans_30_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_30_shiftAmt_T_2 = ans_30_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_30_shiftAmt = ans_30_expRaw > 6'h3 ? _ans_30_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_30_mantissaRaw_T = ans_30_absClipped >> ans_30_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_30_mantissaRaw = _ans_30_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_30_mantissa = ans_30_expRaw >= 6'h3 ? ans_30_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_30_expAdjusted = ans_30_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_30_exp_T_4 = ans_30_expAdjusted > 7'hf ? 4'hf : ans_30_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_30_exp = ans_30_isZero ? 4'h0 : _ans_30_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_30_fp8 = {ans_30_clippedX[31],ans_30_exp,ans_30_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_31 = {24'h0,linear_bias_31}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_31 = tempSum_31 + biasExtended_31; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_31_sign = sum32_31[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_31_absX_T = ~sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_31_absX_T_2 = _ans_31_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_31_absX = ans_31_sign ? _ans_31_absX_T_2 : sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_31_shiftedX_T_1 = _GEN_10432 - ans_31_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_31_shiftedX_T_3 = ans_31_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_31_shiftedX = ans_31_sign ? _ans_31_shiftedX_T_1 : _ans_31_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_31_scaledX_T_1 = ans_31_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_31_scaledX = _ans_31_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_31_clippedX_T_2 = ans_31_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_31_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_31_clippedX = ans_31_scaledX > 49'h1c0 ? 49'h1c0 : _ans_31_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_31_absClipped_T_1 = ~ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_31_absClipped_T_3 = _ans_31_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_31_absClipped = ans_31_clippedX[31] ? _ans_31_absClipped_T_3 : ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_31_isZero = ans_31_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10775 = {{16'd0}, ans_31_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_4 = _GEN_10775 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_6 = {ans_31_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_8 = _ans_31_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_9 = _ans_31_leadingZeros_T_4 | _ans_31_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10776 = {{8'd0}, _ans_31_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_14 = _GEN_10776 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_16 = {_ans_31_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_18 = _ans_31_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_19 = _ans_31_leadingZeros_T_14 | _ans_31_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10777 = {{4'd0}, _ans_31_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_24 = _GEN_10777 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_26 = {_ans_31_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_28 = _ans_31_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_29 = _ans_31_leadingZeros_T_24 | _ans_31_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10778 = {{2'd0}, _ans_31_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_34 = _GEN_10778 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_36 = {_ans_31_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_38 = _ans_31_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_39 = _ans_31_leadingZeros_T_34 | _ans_31_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10779 = {{1'd0}, _ans_31_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_44 = _GEN_10779 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_46 = {_ans_31_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_48 = _ans_31_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_31_leadingZeros_T_49 = _ans_31_leadingZeros_T_44 | _ans_31_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10780 = {{8'd0}, ans_31_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_55 = _GEN_10780 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_57 = {ans_31_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_59 = _ans_31_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_60 = _ans_31_leadingZeros_T_55 | _ans_31_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10781 = {{4'd0}, _ans_31_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_65 = _GEN_10781 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_67 = {_ans_31_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_69 = _ans_31_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_70 = _ans_31_leadingZeros_T_65 | _ans_31_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10782 = {{2'd0}, _ans_31_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_75 = _GEN_10782 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_77 = {_ans_31_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_79 = _ans_31_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_80 = _ans_31_leadingZeros_T_75 | _ans_31_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10783 = {{1'd0}, _ans_31_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_85 = _GEN_10783 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_87 = {_ans_31_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_89 = _ans_31_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_31_leadingZeros_T_90 = _ans_31_leadingZeros_T_85 | _ans_31_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_31_leadingZeros_T_93 = {_ans_31_leadingZeros_T_49,_ans_31_leadingZeros_T_90,ans_31_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_31_leadingZeros_T_143 = _ans_31_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_144 = _ans_31_leadingZeros_T_93[46] ? 6'h2e : _ans_31_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_145 = _ans_31_leadingZeros_T_93[45] ? 6'h2d : _ans_31_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_146 = _ans_31_leadingZeros_T_93[44] ? 6'h2c : _ans_31_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_147 = _ans_31_leadingZeros_T_93[43] ? 6'h2b : _ans_31_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_148 = _ans_31_leadingZeros_T_93[42] ? 6'h2a : _ans_31_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_149 = _ans_31_leadingZeros_T_93[41] ? 6'h29 : _ans_31_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_150 = _ans_31_leadingZeros_T_93[40] ? 6'h28 : _ans_31_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_151 = _ans_31_leadingZeros_T_93[39] ? 6'h27 : _ans_31_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_152 = _ans_31_leadingZeros_T_93[38] ? 6'h26 : _ans_31_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_153 = _ans_31_leadingZeros_T_93[37] ? 6'h25 : _ans_31_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_154 = _ans_31_leadingZeros_T_93[36] ? 6'h24 : _ans_31_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_155 = _ans_31_leadingZeros_T_93[35] ? 6'h23 : _ans_31_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_156 = _ans_31_leadingZeros_T_93[34] ? 6'h22 : _ans_31_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_157 = _ans_31_leadingZeros_T_93[33] ? 6'h21 : _ans_31_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_158 = _ans_31_leadingZeros_T_93[32] ? 6'h20 : _ans_31_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_159 = _ans_31_leadingZeros_T_93[31] ? 6'h1f : _ans_31_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_160 = _ans_31_leadingZeros_T_93[30] ? 6'h1e : _ans_31_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_161 = _ans_31_leadingZeros_T_93[29] ? 6'h1d : _ans_31_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_162 = _ans_31_leadingZeros_T_93[28] ? 6'h1c : _ans_31_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_163 = _ans_31_leadingZeros_T_93[27] ? 6'h1b : _ans_31_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_164 = _ans_31_leadingZeros_T_93[26] ? 6'h1a : _ans_31_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_165 = _ans_31_leadingZeros_T_93[25] ? 6'h19 : _ans_31_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_166 = _ans_31_leadingZeros_T_93[24] ? 6'h18 : _ans_31_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_167 = _ans_31_leadingZeros_T_93[23] ? 6'h17 : _ans_31_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_168 = _ans_31_leadingZeros_T_93[22] ? 6'h16 : _ans_31_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_169 = _ans_31_leadingZeros_T_93[21] ? 6'h15 : _ans_31_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_170 = _ans_31_leadingZeros_T_93[20] ? 6'h14 : _ans_31_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_171 = _ans_31_leadingZeros_T_93[19] ? 6'h13 : _ans_31_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_172 = _ans_31_leadingZeros_T_93[18] ? 6'h12 : _ans_31_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_173 = _ans_31_leadingZeros_T_93[17] ? 6'h11 : _ans_31_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_174 = _ans_31_leadingZeros_T_93[16] ? 6'h10 : _ans_31_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_175 = _ans_31_leadingZeros_T_93[15] ? 6'hf : _ans_31_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_176 = _ans_31_leadingZeros_T_93[14] ? 6'he : _ans_31_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_177 = _ans_31_leadingZeros_T_93[13] ? 6'hd : _ans_31_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_178 = _ans_31_leadingZeros_T_93[12] ? 6'hc : _ans_31_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_179 = _ans_31_leadingZeros_T_93[11] ? 6'hb : _ans_31_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_180 = _ans_31_leadingZeros_T_93[10] ? 6'ha : _ans_31_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_181 = _ans_31_leadingZeros_T_93[9] ? 6'h9 : _ans_31_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_182 = _ans_31_leadingZeros_T_93[8] ? 6'h8 : _ans_31_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_183 = _ans_31_leadingZeros_T_93[7] ? 6'h7 : _ans_31_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_184 = _ans_31_leadingZeros_T_93[6] ? 6'h6 : _ans_31_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_185 = _ans_31_leadingZeros_T_93[5] ? 6'h5 : _ans_31_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_186 = _ans_31_leadingZeros_T_93[4] ? 6'h4 : _ans_31_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_187 = _ans_31_leadingZeros_T_93[3] ? 6'h3 : _ans_31_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_188 = _ans_31_leadingZeros_T_93[2] ? 6'h2 : _ans_31_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_189 = _ans_31_leadingZeros_T_93[1] ? 6'h1 : _ans_31_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_31_leadingZeros = _ans_31_leadingZeros_T_93[0] ? 6'h0 : _ans_31_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_expRaw_T_1 = 6'h1f - ans_31_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_31_expRaw = ans_31_isZero ? 6'h0 : _ans_31_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_31_shiftAmt_T_2 = ans_31_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_31_shiftAmt = ans_31_expRaw > 6'h3 ? _ans_31_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_31_mantissaRaw_T = ans_31_absClipped >> ans_31_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_31_mantissaRaw = _ans_31_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_31_mantissa = ans_31_expRaw >= 6'h3 ? ans_31_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_31_expAdjusted = ans_31_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_31_exp_T_4 = ans_31_expAdjusted > 7'hf ? 4'hf : ans_31_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_31_exp = ans_31_isZero ? 4'h0 : _ans_31_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_31_fp8 = {ans_31_clippedX[31],ans_31_exp,ans_31_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_32 = {24'h0,linear_bias_32}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_32 = tempSum_32 + biasExtended_32; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_32_sign = sum32_32[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_32_absX_T = ~sum32_32; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_32_absX_T_2 = _ans_32_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_32_absX = ans_32_sign ? _ans_32_absX_T_2 : sum32_32; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_32_shiftedX_T_1 = _GEN_10432 - ans_32_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_32_shiftedX_T_3 = ans_32_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_32_shiftedX = ans_32_sign ? _ans_32_shiftedX_T_1 : _ans_32_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_32_scaledX_T_1 = ans_32_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_32_scaledX = _ans_32_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_32_clippedX_T_2 = ans_32_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_32_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_32_clippedX = ans_32_scaledX > 49'h1c0 ? 49'h1c0 : _ans_32_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_32_absClipped_T_1 = ~ans_32_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_32_absClipped_T_3 = _ans_32_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_32_absClipped = ans_32_clippedX[31] ? _ans_32_absClipped_T_3 : ans_32_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_32_isZero = ans_32_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10786 = {{16'd0}, ans_32_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_4 = _GEN_10786 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_6 = {ans_32_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_8 = _ans_32_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_9 = _ans_32_leadingZeros_T_4 | _ans_32_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10787 = {{8'd0}, _ans_32_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_14 = _GEN_10787 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_16 = {_ans_32_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_18 = _ans_32_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_19 = _ans_32_leadingZeros_T_14 | _ans_32_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10788 = {{4'd0}, _ans_32_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_24 = _GEN_10788 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_26 = {_ans_32_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_28 = _ans_32_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_29 = _ans_32_leadingZeros_T_24 | _ans_32_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10789 = {{2'd0}, _ans_32_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_34 = _GEN_10789 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_36 = {_ans_32_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_38 = _ans_32_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_39 = _ans_32_leadingZeros_T_34 | _ans_32_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10790 = {{1'd0}, _ans_32_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_44 = _GEN_10790 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_46 = {_ans_32_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_48 = _ans_32_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_32_leadingZeros_T_49 = _ans_32_leadingZeros_T_44 | _ans_32_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10791 = {{8'd0}, ans_32_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_55 = _GEN_10791 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_57 = {ans_32_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_59 = _ans_32_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_60 = _ans_32_leadingZeros_T_55 | _ans_32_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10792 = {{4'd0}, _ans_32_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_65 = _GEN_10792 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_67 = {_ans_32_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_69 = _ans_32_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_70 = _ans_32_leadingZeros_T_65 | _ans_32_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10793 = {{2'd0}, _ans_32_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_75 = _GEN_10793 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_77 = {_ans_32_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_79 = _ans_32_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_80 = _ans_32_leadingZeros_T_75 | _ans_32_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10794 = {{1'd0}, _ans_32_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_85 = _GEN_10794 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_87 = {_ans_32_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_89 = _ans_32_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_32_leadingZeros_T_90 = _ans_32_leadingZeros_T_85 | _ans_32_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_32_leadingZeros_T_93 = {_ans_32_leadingZeros_T_49,_ans_32_leadingZeros_T_90,ans_32_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_32_leadingZeros_T_143 = _ans_32_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_144 = _ans_32_leadingZeros_T_93[46] ? 6'h2e : _ans_32_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_145 = _ans_32_leadingZeros_T_93[45] ? 6'h2d : _ans_32_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_146 = _ans_32_leadingZeros_T_93[44] ? 6'h2c : _ans_32_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_147 = _ans_32_leadingZeros_T_93[43] ? 6'h2b : _ans_32_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_148 = _ans_32_leadingZeros_T_93[42] ? 6'h2a : _ans_32_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_149 = _ans_32_leadingZeros_T_93[41] ? 6'h29 : _ans_32_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_150 = _ans_32_leadingZeros_T_93[40] ? 6'h28 : _ans_32_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_151 = _ans_32_leadingZeros_T_93[39] ? 6'h27 : _ans_32_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_152 = _ans_32_leadingZeros_T_93[38] ? 6'h26 : _ans_32_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_153 = _ans_32_leadingZeros_T_93[37] ? 6'h25 : _ans_32_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_154 = _ans_32_leadingZeros_T_93[36] ? 6'h24 : _ans_32_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_155 = _ans_32_leadingZeros_T_93[35] ? 6'h23 : _ans_32_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_156 = _ans_32_leadingZeros_T_93[34] ? 6'h22 : _ans_32_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_157 = _ans_32_leadingZeros_T_93[33] ? 6'h21 : _ans_32_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_158 = _ans_32_leadingZeros_T_93[32] ? 6'h20 : _ans_32_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_159 = _ans_32_leadingZeros_T_93[31] ? 6'h1f : _ans_32_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_160 = _ans_32_leadingZeros_T_93[30] ? 6'h1e : _ans_32_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_161 = _ans_32_leadingZeros_T_93[29] ? 6'h1d : _ans_32_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_162 = _ans_32_leadingZeros_T_93[28] ? 6'h1c : _ans_32_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_163 = _ans_32_leadingZeros_T_93[27] ? 6'h1b : _ans_32_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_164 = _ans_32_leadingZeros_T_93[26] ? 6'h1a : _ans_32_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_165 = _ans_32_leadingZeros_T_93[25] ? 6'h19 : _ans_32_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_166 = _ans_32_leadingZeros_T_93[24] ? 6'h18 : _ans_32_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_167 = _ans_32_leadingZeros_T_93[23] ? 6'h17 : _ans_32_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_168 = _ans_32_leadingZeros_T_93[22] ? 6'h16 : _ans_32_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_169 = _ans_32_leadingZeros_T_93[21] ? 6'h15 : _ans_32_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_170 = _ans_32_leadingZeros_T_93[20] ? 6'h14 : _ans_32_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_171 = _ans_32_leadingZeros_T_93[19] ? 6'h13 : _ans_32_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_172 = _ans_32_leadingZeros_T_93[18] ? 6'h12 : _ans_32_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_173 = _ans_32_leadingZeros_T_93[17] ? 6'h11 : _ans_32_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_174 = _ans_32_leadingZeros_T_93[16] ? 6'h10 : _ans_32_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_175 = _ans_32_leadingZeros_T_93[15] ? 6'hf : _ans_32_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_176 = _ans_32_leadingZeros_T_93[14] ? 6'he : _ans_32_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_177 = _ans_32_leadingZeros_T_93[13] ? 6'hd : _ans_32_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_178 = _ans_32_leadingZeros_T_93[12] ? 6'hc : _ans_32_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_179 = _ans_32_leadingZeros_T_93[11] ? 6'hb : _ans_32_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_180 = _ans_32_leadingZeros_T_93[10] ? 6'ha : _ans_32_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_181 = _ans_32_leadingZeros_T_93[9] ? 6'h9 : _ans_32_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_182 = _ans_32_leadingZeros_T_93[8] ? 6'h8 : _ans_32_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_183 = _ans_32_leadingZeros_T_93[7] ? 6'h7 : _ans_32_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_184 = _ans_32_leadingZeros_T_93[6] ? 6'h6 : _ans_32_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_185 = _ans_32_leadingZeros_T_93[5] ? 6'h5 : _ans_32_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_186 = _ans_32_leadingZeros_T_93[4] ? 6'h4 : _ans_32_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_187 = _ans_32_leadingZeros_T_93[3] ? 6'h3 : _ans_32_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_188 = _ans_32_leadingZeros_T_93[2] ? 6'h2 : _ans_32_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_leadingZeros_T_189 = _ans_32_leadingZeros_T_93[1] ? 6'h1 : _ans_32_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_32_leadingZeros = _ans_32_leadingZeros_T_93[0] ? 6'h0 : _ans_32_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_32_expRaw_T_1 = 6'h1f - ans_32_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_32_expRaw = ans_32_isZero ? 6'h0 : _ans_32_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_32_shiftAmt_T_2 = ans_32_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_32_shiftAmt = ans_32_expRaw > 6'h3 ? _ans_32_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_32_mantissaRaw_T = ans_32_absClipped >> ans_32_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_32_mantissaRaw = _ans_32_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_32_mantissa = ans_32_expRaw >= 6'h3 ? ans_32_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_32_expAdjusted = ans_32_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_32_exp_T_4 = ans_32_expAdjusted > 7'hf ? 4'hf : ans_32_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_32_exp = ans_32_isZero ? 4'h0 : _ans_32_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_32_fp8 = {ans_32_clippedX[31],ans_32_exp,ans_32_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_33 = {24'h0,linear_bias_33}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_33 = tempSum_33 + biasExtended_33; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_33_sign = sum32_33[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_33_absX_T = ~sum32_33; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_33_absX_T_2 = _ans_33_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_33_absX = ans_33_sign ? _ans_33_absX_T_2 : sum32_33; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_33_shiftedX_T_1 = _GEN_10432 - ans_33_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_33_shiftedX_T_3 = ans_33_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_33_shiftedX = ans_33_sign ? _ans_33_shiftedX_T_1 : _ans_33_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_33_scaledX_T_1 = ans_33_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_33_scaledX = _ans_33_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_33_clippedX_T_2 = ans_33_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_33_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_33_clippedX = ans_33_scaledX > 49'h1c0 ? 49'h1c0 : _ans_33_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_33_absClipped_T_1 = ~ans_33_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_33_absClipped_T_3 = _ans_33_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_33_absClipped = ans_33_clippedX[31] ? _ans_33_absClipped_T_3 : ans_33_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_33_isZero = ans_33_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10797 = {{16'd0}, ans_33_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_4 = _GEN_10797 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_6 = {ans_33_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_8 = _ans_33_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_9 = _ans_33_leadingZeros_T_4 | _ans_33_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10798 = {{8'd0}, _ans_33_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_14 = _GEN_10798 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_16 = {_ans_33_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_18 = _ans_33_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_19 = _ans_33_leadingZeros_T_14 | _ans_33_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10799 = {{4'd0}, _ans_33_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_24 = _GEN_10799 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_26 = {_ans_33_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_28 = _ans_33_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_29 = _ans_33_leadingZeros_T_24 | _ans_33_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10800 = {{2'd0}, _ans_33_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_34 = _GEN_10800 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_36 = {_ans_33_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_38 = _ans_33_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_39 = _ans_33_leadingZeros_T_34 | _ans_33_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10801 = {{1'd0}, _ans_33_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_44 = _GEN_10801 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_46 = {_ans_33_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_48 = _ans_33_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_33_leadingZeros_T_49 = _ans_33_leadingZeros_T_44 | _ans_33_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10802 = {{8'd0}, ans_33_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_55 = _GEN_10802 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_57 = {ans_33_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_59 = _ans_33_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_60 = _ans_33_leadingZeros_T_55 | _ans_33_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10803 = {{4'd0}, _ans_33_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_65 = _GEN_10803 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_67 = {_ans_33_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_69 = _ans_33_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_70 = _ans_33_leadingZeros_T_65 | _ans_33_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10804 = {{2'd0}, _ans_33_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_75 = _GEN_10804 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_77 = {_ans_33_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_79 = _ans_33_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_80 = _ans_33_leadingZeros_T_75 | _ans_33_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10805 = {{1'd0}, _ans_33_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_85 = _GEN_10805 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_87 = {_ans_33_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_89 = _ans_33_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_33_leadingZeros_T_90 = _ans_33_leadingZeros_T_85 | _ans_33_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_33_leadingZeros_T_93 = {_ans_33_leadingZeros_T_49,_ans_33_leadingZeros_T_90,ans_33_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_33_leadingZeros_T_143 = _ans_33_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_144 = _ans_33_leadingZeros_T_93[46] ? 6'h2e : _ans_33_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_145 = _ans_33_leadingZeros_T_93[45] ? 6'h2d : _ans_33_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_146 = _ans_33_leadingZeros_T_93[44] ? 6'h2c : _ans_33_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_147 = _ans_33_leadingZeros_T_93[43] ? 6'h2b : _ans_33_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_148 = _ans_33_leadingZeros_T_93[42] ? 6'h2a : _ans_33_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_149 = _ans_33_leadingZeros_T_93[41] ? 6'h29 : _ans_33_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_150 = _ans_33_leadingZeros_T_93[40] ? 6'h28 : _ans_33_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_151 = _ans_33_leadingZeros_T_93[39] ? 6'h27 : _ans_33_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_152 = _ans_33_leadingZeros_T_93[38] ? 6'h26 : _ans_33_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_153 = _ans_33_leadingZeros_T_93[37] ? 6'h25 : _ans_33_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_154 = _ans_33_leadingZeros_T_93[36] ? 6'h24 : _ans_33_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_155 = _ans_33_leadingZeros_T_93[35] ? 6'h23 : _ans_33_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_156 = _ans_33_leadingZeros_T_93[34] ? 6'h22 : _ans_33_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_157 = _ans_33_leadingZeros_T_93[33] ? 6'h21 : _ans_33_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_158 = _ans_33_leadingZeros_T_93[32] ? 6'h20 : _ans_33_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_159 = _ans_33_leadingZeros_T_93[31] ? 6'h1f : _ans_33_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_160 = _ans_33_leadingZeros_T_93[30] ? 6'h1e : _ans_33_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_161 = _ans_33_leadingZeros_T_93[29] ? 6'h1d : _ans_33_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_162 = _ans_33_leadingZeros_T_93[28] ? 6'h1c : _ans_33_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_163 = _ans_33_leadingZeros_T_93[27] ? 6'h1b : _ans_33_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_164 = _ans_33_leadingZeros_T_93[26] ? 6'h1a : _ans_33_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_165 = _ans_33_leadingZeros_T_93[25] ? 6'h19 : _ans_33_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_166 = _ans_33_leadingZeros_T_93[24] ? 6'h18 : _ans_33_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_167 = _ans_33_leadingZeros_T_93[23] ? 6'h17 : _ans_33_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_168 = _ans_33_leadingZeros_T_93[22] ? 6'h16 : _ans_33_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_169 = _ans_33_leadingZeros_T_93[21] ? 6'h15 : _ans_33_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_170 = _ans_33_leadingZeros_T_93[20] ? 6'h14 : _ans_33_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_171 = _ans_33_leadingZeros_T_93[19] ? 6'h13 : _ans_33_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_172 = _ans_33_leadingZeros_T_93[18] ? 6'h12 : _ans_33_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_173 = _ans_33_leadingZeros_T_93[17] ? 6'h11 : _ans_33_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_174 = _ans_33_leadingZeros_T_93[16] ? 6'h10 : _ans_33_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_175 = _ans_33_leadingZeros_T_93[15] ? 6'hf : _ans_33_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_176 = _ans_33_leadingZeros_T_93[14] ? 6'he : _ans_33_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_177 = _ans_33_leadingZeros_T_93[13] ? 6'hd : _ans_33_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_178 = _ans_33_leadingZeros_T_93[12] ? 6'hc : _ans_33_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_179 = _ans_33_leadingZeros_T_93[11] ? 6'hb : _ans_33_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_180 = _ans_33_leadingZeros_T_93[10] ? 6'ha : _ans_33_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_181 = _ans_33_leadingZeros_T_93[9] ? 6'h9 : _ans_33_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_182 = _ans_33_leadingZeros_T_93[8] ? 6'h8 : _ans_33_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_183 = _ans_33_leadingZeros_T_93[7] ? 6'h7 : _ans_33_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_184 = _ans_33_leadingZeros_T_93[6] ? 6'h6 : _ans_33_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_185 = _ans_33_leadingZeros_T_93[5] ? 6'h5 : _ans_33_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_186 = _ans_33_leadingZeros_T_93[4] ? 6'h4 : _ans_33_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_187 = _ans_33_leadingZeros_T_93[3] ? 6'h3 : _ans_33_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_188 = _ans_33_leadingZeros_T_93[2] ? 6'h2 : _ans_33_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_leadingZeros_T_189 = _ans_33_leadingZeros_T_93[1] ? 6'h1 : _ans_33_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_33_leadingZeros = _ans_33_leadingZeros_T_93[0] ? 6'h0 : _ans_33_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_33_expRaw_T_1 = 6'h1f - ans_33_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_33_expRaw = ans_33_isZero ? 6'h0 : _ans_33_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_33_shiftAmt_T_2 = ans_33_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_33_shiftAmt = ans_33_expRaw > 6'h3 ? _ans_33_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_33_mantissaRaw_T = ans_33_absClipped >> ans_33_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_33_mantissaRaw = _ans_33_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_33_mantissa = ans_33_expRaw >= 6'h3 ? ans_33_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_33_expAdjusted = ans_33_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_33_exp_T_4 = ans_33_expAdjusted > 7'hf ? 4'hf : ans_33_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_33_exp = ans_33_isZero ? 4'h0 : _ans_33_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_33_fp8 = {ans_33_clippedX[31],ans_33_exp,ans_33_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_34 = {24'h0,linear_bias_34}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_34 = tempSum_34 + biasExtended_34; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_34_sign = sum32_34[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_34_absX_T = ~sum32_34; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_34_absX_T_2 = _ans_34_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_34_absX = ans_34_sign ? _ans_34_absX_T_2 : sum32_34; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_34_shiftedX_T_1 = _GEN_10432 - ans_34_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_34_shiftedX_T_3 = ans_34_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_34_shiftedX = ans_34_sign ? _ans_34_shiftedX_T_1 : _ans_34_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_34_scaledX_T_1 = ans_34_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_34_scaledX = _ans_34_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_34_clippedX_T_2 = ans_34_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_34_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_34_clippedX = ans_34_scaledX > 49'h1c0 ? 49'h1c0 : _ans_34_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_34_absClipped_T_1 = ~ans_34_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_34_absClipped_T_3 = _ans_34_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_34_absClipped = ans_34_clippedX[31] ? _ans_34_absClipped_T_3 : ans_34_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_34_isZero = ans_34_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10808 = {{16'd0}, ans_34_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_4 = _GEN_10808 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_6 = {ans_34_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_8 = _ans_34_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_9 = _ans_34_leadingZeros_T_4 | _ans_34_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10809 = {{8'd0}, _ans_34_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_14 = _GEN_10809 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_16 = {_ans_34_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_18 = _ans_34_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_19 = _ans_34_leadingZeros_T_14 | _ans_34_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10810 = {{4'd0}, _ans_34_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_24 = _GEN_10810 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_26 = {_ans_34_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_28 = _ans_34_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_29 = _ans_34_leadingZeros_T_24 | _ans_34_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10811 = {{2'd0}, _ans_34_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_34 = _GEN_10811 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_36 = {_ans_34_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_38 = _ans_34_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_39 = _ans_34_leadingZeros_T_34 | _ans_34_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10812 = {{1'd0}, _ans_34_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_44 = _GEN_10812 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_46 = {_ans_34_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_48 = _ans_34_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_34_leadingZeros_T_49 = _ans_34_leadingZeros_T_44 | _ans_34_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10813 = {{8'd0}, ans_34_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_55 = _GEN_10813 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_57 = {ans_34_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_59 = _ans_34_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_60 = _ans_34_leadingZeros_T_55 | _ans_34_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10814 = {{4'd0}, _ans_34_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_65 = _GEN_10814 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_67 = {_ans_34_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_69 = _ans_34_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_70 = _ans_34_leadingZeros_T_65 | _ans_34_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10815 = {{2'd0}, _ans_34_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_75 = _GEN_10815 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_77 = {_ans_34_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_79 = _ans_34_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_80 = _ans_34_leadingZeros_T_75 | _ans_34_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10816 = {{1'd0}, _ans_34_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_85 = _GEN_10816 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_87 = {_ans_34_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_89 = _ans_34_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_34_leadingZeros_T_90 = _ans_34_leadingZeros_T_85 | _ans_34_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_34_leadingZeros_T_93 = {_ans_34_leadingZeros_T_49,_ans_34_leadingZeros_T_90,ans_34_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_34_leadingZeros_T_143 = _ans_34_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_144 = _ans_34_leadingZeros_T_93[46] ? 6'h2e : _ans_34_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_145 = _ans_34_leadingZeros_T_93[45] ? 6'h2d : _ans_34_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_146 = _ans_34_leadingZeros_T_93[44] ? 6'h2c : _ans_34_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_147 = _ans_34_leadingZeros_T_93[43] ? 6'h2b : _ans_34_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_148 = _ans_34_leadingZeros_T_93[42] ? 6'h2a : _ans_34_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_149 = _ans_34_leadingZeros_T_93[41] ? 6'h29 : _ans_34_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_150 = _ans_34_leadingZeros_T_93[40] ? 6'h28 : _ans_34_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_151 = _ans_34_leadingZeros_T_93[39] ? 6'h27 : _ans_34_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_152 = _ans_34_leadingZeros_T_93[38] ? 6'h26 : _ans_34_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_153 = _ans_34_leadingZeros_T_93[37] ? 6'h25 : _ans_34_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_154 = _ans_34_leadingZeros_T_93[36] ? 6'h24 : _ans_34_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_155 = _ans_34_leadingZeros_T_93[35] ? 6'h23 : _ans_34_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_156 = _ans_34_leadingZeros_T_93[34] ? 6'h22 : _ans_34_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_157 = _ans_34_leadingZeros_T_93[33] ? 6'h21 : _ans_34_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_158 = _ans_34_leadingZeros_T_93[32] ? 6'h20 : _ans_34_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_159 = _ans_34_leadingZeros_T_93[31] ? 6'h1f : _ans_34_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_160 = _ans_34_leadingZeros_T_93[30] ? 6'h1e : _ans_34_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_161 = _ans_34_leadingZeros_T_93[29] ? 6'h1d : _ans_34_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_162 = _ans_34_leadingZeros_T_93[28] ? 6'h1c : _ans_34_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_163 = _ans_34_leadingZeros_T_93[27] ? 6'h1b : _ans_34_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_164 = _ans_34_leadingZeros_T_93[26] ? 6'h1a : _ans_34_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_165 = _ans_34_leadingZeros_T_93[25] ? 6'h19 : _ans_34_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_166 = _ans_34_leadingZeros_T_93[24] ? 6'h18 : _ans_34_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_167 = _ans_34_leadingZeros_T_93[23] ? 6'h17 : _ans_34_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_168 = _ans_34_leadingZeros_T_93[22] ? 6'h16 : _ans_34_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_169 = _ans_34_leadingZeros_T_93[21] ? 6'h15 : _ans_34_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_170 = _ans_34_leadingZeros_T_93[20] ? 6'h14 : _ans_34_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_171 = _ans_34_leadingZeros_T_93[19] ? 6'h13 : _ans_34_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_172 = _ans_34_leadingZeros_T_93[18] ? 6'h12 : _ans_34_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_173 = _ans_34_leadingZeros_T_93[17] ? 6'h11 : _ans_34_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_174 = _ans_34_leadingZeros_T_93[16] ? 6'h10 : _ans_34_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_175 = _ans_34_leadingZeros_T_93[15] ? 6'hf : _ans_34_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_176 = _ans_34_leadingZeros_T_93[14] ? 6'he : _ans_34_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_177 = _ans_34_leadingZeros_T_93[13] ? 6'hd : _ans_34_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_178 = _ans_34_leadingZeros_T_93[12] ? 6'hc : _ans_34_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_179 = _ans_34_leadingZeros_T_93[11] ? 6'hb : _ans_34_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_180 = _ans_34_leadingZeros_T_93[10] ? 6'ha : _ans_34_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_181 = _ans_34_leadingZeros_T_93[9] ? 6'h9 : _ans_34_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_182 = _ans_34_leadingZeros_T_93[8] ? 6'h8 : _ans_34_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_183 = _ans_34_leadingZeros_T_93[7] ? 6'h7 : _ans_34_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_184 = _ans_34_leadingZeros_T_93[6] ? 6'h6 : _ans_34_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_185 = _ans_34_leadingZeros_T_93[5] ? 6'h5 : _ans_34_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_186 = _ans_34_leadingZeros_T_93[4] ? 6'h4 : _ans_34_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_187 = _ans_34_leadingZeros_T_93[3] ? 6'h3 : _ans_34_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_188 = _ans_34_leadingZeros_T_93[2] ? 6'h2 : _ans_34_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_leadingZeros_T_189 = _ans_34_leadingZeros_T_93[1] ? 6'h1 : _ans_34_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_34_leadingZeros = _ans_34_leadingZeros_T_93[0] ? 6'h0 : _ans_34_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_34_expRaw_T_1 = 6'h1f - ans_34_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_34_expRaw = ans_34_isZero ? 6'h0 : _ans_34_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_34_shiftAmt_T_2 = ans_34_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_34_shiftAmt = ans_34_expRaw > 6'h3 ? _ans_34_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_34_mantissaRaw_T = ans_34_absClipped >> ans_34_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_34_mantissaRaw = _ans_34_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_34_mantissa = ans_34_expRaw >= 6'h3 ? ans_34_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_34_expAdjusted = ans_34_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_34_exp_T_4 = ans_34_expAdjusted > 7'hf ? 4'hf : ans_34_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_34_exp = ans_34_isZero ? 4'h0 : _ans_34_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_34_fp8 = {ans_34_clippedX[31],ans_34_exp,ans_34_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_35 = {24'h0,linear_bias_35}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_35 = tempSum_35 + biasExtended_35; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_35_sign = sum32_35[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_35_absX_T = ~sum32_35; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_35_absX_T_2 = _ans_35_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_35_absX = ans_35_sign ? _ans_35_absX_T_2 : sum32_35; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_35_shiftedX_T_1 = _GEN_10432 - ans_35_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_35_shiftedX_T_3 = ans_35_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_35_shiftedX = ans_35_sign ? _ans_35_shiftedX_T_1 : _ans_35_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_35_scaledX_T_1 = ans_35_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_35_scaledX = _ans_35_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_35_clippedX_T_2 = ans_35_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_35_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_35_clippedX = ans_35_scaledX > 49'h1c0 ? 49'h1c0 : _ans_35_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_35_absClipped_T_1 = ~ans_35_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_35_absClipped_T_3 = _ans_35_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_35_absClipped = ans_35_clippedX[31] ? _ans_35_absClipped_T_3 : ans_35_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_35_isZero = ans_35_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10819 = {{16'd0}, ans_35_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_4 = _GEN_10819 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_6 = {ans_35_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_8 = _ans_35_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_9 = _ans_35_leadingZeros_T_4 | _ans_35_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10820 = {{8'd0}, _ans_35_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_14 = _GEN_10820 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_16 = {_ans_35_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_18 = _ans_35_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_19 = _ans_35_leadingZeros_T_14 | _ans_35_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10821 = {{4'd0}, _ans_35_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_24 = _GEN_10821 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_26 = {_ans_35_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_28 = _ans_35_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_29 = _ans_35_leadingZeros_T_24 | _ans_35_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10822 = {{2'd0}, _ans_35_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_34 = _GEN_10822 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_36 = {_ans_35_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_38 = _ans_35_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_39 = _ans_35_leadingZeros_T_34 | _ans_35_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10823 = {{1'd0}, _ans_35_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_44 = _GEN_10823 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_46 = {_ans_35_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_48 = _ans_35_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_35_leadingZeros_T_49 = _ans_35_leadingZeros_T_44 | _ans_35_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10824 = {{8'd0}, ans_35_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_55 = _GEN_10824 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_57 = {ans_35_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_59 = _ans_35_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_60 = _ans_35_leadingZeros_T_55 | _ans_35_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10825 = {{4'd0}, _ans_35_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_65 = _GEN_10825 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_67 = {_ans_35_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_69 = _ans_35_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_70 = _ans_35_leadingZeros_T_65 | _ans_35_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10826 = {{2'd0}, _ans_35_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_75 = _GEN_10826 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_77 = {_ans_35_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_79 = _ans_35_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_80 = _ans_35_leadingZeros_T_75 | _ans_35_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10827 = {{1'd0}, _ans_35_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_85 = _GEN_10827 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_87 = {_ans_35_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_89 = _ans_35_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_35_leadingZeros_T_90 = _ans_35_leadingZeros_T_85 | _ans_35_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_35_leadingZeros_T_93 = {_ans_35_leadingZeros_T_49,_ans_35_leadingZeros_T_90,ans_35_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_35_leadingZeros_T_143 = _ans_35_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_144 = _ans_35_leadingZeros_T_93[46] ? 6'h2e : _ans_35_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_145 = _ans_35_leadingZeros_T_93[45] ? 6'h2d : _ans_35_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_146 = _ans_35_leadingZeros_T_93[44] ? 6'h2c : _ans_35_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_147 = _ans_35_leadingZeros_T_93[43] ? 6'h2b : _ans_35_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_148 = _ans_35_leadingZeros_T_93[42] ? 6'h2a : _ans_35_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_149 = _ans_35_leadingZeros_T_93[41] ? 6'h29 : _ans_35_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_150 = _ans_35_leadingZeros_T_93[40] ? 6'h28 : _ans_35_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_151 = _ans_35_leadingZeros_T_93[39] ? 6'h27 : _ans_35_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_152 = _ans_35_leadingZeros_T_93[38] ? 6'h26 : _ans_35_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_153 = _ans_35_leadingZeros_T_93[37] ? 6'h25 : _ans_35_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_154 = _ans_35_leadingZeros_T_93[36] ? 6'h24 : _ans_35_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_155 = _ans_35_leadingZeros_T_93[35] ? 6'h23 : _ans_35_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_156 = _ans_35_leadingZeros_T_93[34] ? 6'h22 : _ans_35_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_157 = _ans_35_leadingZeros_T_93[33] ? 6'h21 : _ans_35_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_158 = _ans_35_leadingZeros_T_93[32] ? 6'h20 : _ans_35_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_159 = _ans_35_leadingZeros_T_93[31] ? 6'h1f : _ans_35_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_160 = _ans_35_leadingZeros_T_93[30] ? 6'h1e : _ans_35_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_161 = _ans_35_leadingZeros_T_93[29] ? 6'h1d : _ans_35_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_162 = _ans_35_leadingZeros_T_93[28] ? 6'h1c : _ans_35_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_163 = _ans_35_leadingZeros_T_93[27] ? 6'h1b : _ans_35_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_164 = _ans_35_leadingZeros_T_93[26] ? 6'h1a : _ans_35_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_165 = _ans_35_leadingZeros_T_93[25] ? 6'h19 : _ans_35_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_166 = _ans_35_leadingZeros_T_93[24] ? 6'h18 : _ans_35_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_167 = _ans_35_leadingZeros_T_93[23] ? 6'h17 : _ans_35_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_168 = _ans_35_leadingZeros_T_93[22] ? 6'h16 : _ans_35_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_169 = _ans_35_leadingZeros_T_93[21] ? 6'h15 : _ans_35_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_170 = _ans_35_leadingZeros_T_93[20] ? 6'h14 : _ans_35_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_171 = _ans_35_leadingZeros_T_93[19] ? 6'h13 : _ans_35_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_172 = _ans_35_leadingZeros_T_93[18] ? 6'h12 : _ans_35_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_173 = _ans_35_leadingZeros_T_93[17] ? 6'h11 : _ans_35_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_174 = _ans_35_leadingZeros_T_93[16] ? 6'h10 : _ans_35_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_175 = _ans_35_leadingZeros_T_93[15] ? 6'hf : _ans_35_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_176 = _ans_35_leadingZeros_T_93[14] ? 6'he : _ans_35_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_177 = _ans_35_leadingZeros_T_93[13] ? 6'hd : _ans_35_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_178 = _ans_35_leadingZeros_T_93[12] ? 6'hc : _ans_35_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_179 = _ans_35_leadingZeros_T_93[11] ? 6'hb : _ans_35_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_180 = _ans_35_leadingZeros_T_93[10] ? 6'ha : _ans_35_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_181 = _ans_35_leadingZeros_T_93[9] ? 6'h9 : _ans_35_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_182 = _ans_35_leadingZeros_T_93[8] ? 6'h8 : _ans_35_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_183 = _ans_35_leadingZeros_T_93[7] ? 6'h7 : _ans_35_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_184 = _ans_35_leadingZeros_T_93[6] ? 6'h6 : _ans_35_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_185 = _ans_35_leadingZeros_T_93[5] ? 6'h5 : _ans_35_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_186 = _ans_35_leadingZeros_T_93[4] ? 6'h4 : _ans_35_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_187 = _ans_35_leadingZeros_T_93[3] ? 6'h3 : _ans_35_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_188 = _ans_35_leadingZeros_T_93[2] ? 6'h2 : _ans_35_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_leadingZeros_T_189 = _ans_35_leadingZeros_T_93[1] ? 6'h1 : _ans_35_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_35_leadingZeros = _ans_35_leadingZeros_T_93[0] ? 6'h0 : _ans_35_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_35_expRaw_T_1 = 6'h1f - ans_35_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_35_expRaw = ans_35_isZero ? 6'h0 : _ans_35_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_35_shiftAmt_T_2 = ans_35_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_35_shiftAmt = ans_35_expRaw > 6'h3 ? _ans_35_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_35_mantissaRaw_T = ans_35_absClipped >> ans_35_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_35_mantissaRaw = _ans_35_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_35_mantissa = ans_35_expRaw >= 6'h3 ? ans_35_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_35_expAdjusted = ans_35_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_35_exp_T_4 = ans_35_expAdjusted > 7'hf ? 4'hf : ans_35_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_35_exp = ans_35_isZero ? 4'h0 : _ans_35_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_35_fp8 = {ans_35_clippedX[31],ans_35_exp,ans_35_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_36 = {24'h0,linear_bias_36}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_36 = tempSum_36 + biasExtended_36; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_36_sign = sum32_36[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_36_absX_T = ~sum32_36; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_36_absX_T_2 = _ans_36_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_36_absX = ans_36_sign ? _ans_36_absX_T_2 : sum32_36; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_36_shiftedX_T_1 = _GEN_10432 - ans_36_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_36_shiftedX_T_3 = ans_36_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_36_shiftedX = ans_36_sign ? _ans_36_shiftedX_T_1 : _ans_36_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_36_scaledX_T_1 = ans_36_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_36_scaledX = _ans_36_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_36_clippedX_T_2 = ans_36_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_36_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_36_clippedX = ans_36_scaledX > 49'h1c0 ? 49'h1c0 : _ans_36_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_36_absClipped_T_1 = ~ans_36_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_36_absClipped_T_3 = _ans_36_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_36_absClipped = ans_36_clippedX[31] ? _ans_36_absClipped_T_3 : ans_36_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_36_isZero = ans_36_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10830 = {{16'd0}, ans_36_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_4 = _GEN_10830 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_6 = {ans_36_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_8 = _ans_36_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_9 = _ans_36_leadingZeros_T_4 | _ans_36_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10831 = {{8'd0}, _ans_36_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_14 = _GEN_10831 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_16 = {_ans_36_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_18 = _ans_36_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_19 = _ans_36_leadingZeros_T_14 | _ans_36_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10832 = {{4'd0}, _ans_36_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_24 = _GEN_10832 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_26 = {_ans_36_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_28 = _ans_36_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_29 = _ans_36_leadingZeros_T_24 | _ans_36_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10833 = {{2'd0}, _ans_36_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_34 = _GEN_10833 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_36 = {_ans_36_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_38 = _ans_36_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_39 = _ans_36_leadingZeros_T_34 | _ans_36_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10834 = {{1'd0}, _ans_36_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_44 = _GEN_10834 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_46 = {_ans_36_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_48 = _ans_36_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_36_leadingZeros_T_49 = _ans_36_leadingZeros_T_44 | _ans_36_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10835 = {{8'd0}, ans_36_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_55 = _GEN_10835 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_57 = {ans_36_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_59 = _ans_36_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_60 = _ans_36_leadingZeros_T_55 | _ans_36_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10836 = {{4'd0}, _ans_36_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_65 = _GEN_10836 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_67 = {_ans_36_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_69 = _ans_36_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_70 = _ans_36_leadingZeros_T_65 | _ans_36_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10837 = {{2'd0}, _ans_36_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_75 = _GEN_10837 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_77 = {_ans_36_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_79 = _ans_36_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_80 = _ans_36_leadingZeros_T_75 | _ans_36_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10838 = {{1'd0}, _ans_36_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_85 = _GEN_10838 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_87 = {_ans_36_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_89 = _ans_36_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_36_leadingZeros_T_90 = _ans_36_leadingZeros_T_85 | _ans_36_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_36_leadingZeros_T_93 = {_ans_36_leadingZeros_T_49,_ans_36_leadingZeros_T_90,ans_36_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_36_leadingZeros_T_143 = _ans_36_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_144 = _ans_36_leadingZeros_T_93[46] ? 6'h2e : _ans_36_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_145 = _ans_36_leadingZeros_T_93[45] ? 6'h2d : _ans_36_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_146 = _ans_36_leadingZeros_T_93[44] ? 6'h2c : _ans_36_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_147 = _ans_36_leadingZeros_T_93[43] ? 6'h2b : _ans_36_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_148 = _ans_36_leadingZeros_T_93[42] ? 6'h2a : _ans_36_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_149 = _ans_36_leadingZeros_T_93[41] ? 6'h29 : _ans_36_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_150 = _ans_36_leadingZeros_T_93[40] ? 6'h28 : _ans_36_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_151 = _ans_36_leadingZeros_T_93[39] ? 6'h27 : _ans_36_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_152 = _ans_36_leadingZeros_T_93[38] ? 6'h26 : _ans_36_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_153 = _ans_36_leadingZeros_T_93[37] ? 6'h25 : _ans_36_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_154 = _ans_36_leadingZeros_T_93[36] ? 6'h24 : _ans_36_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_155 = _ans_36_leadingZeros_T_93[35] ? 6'h23 : _ans_36_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_156 = _ans_36_leadingZeros_T_93[34] ? 6'h22 : _ans_36_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_157 = _ans_36_leadingZeros_T_93[33] ? 6'h21 : _ans_36_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_158 = _ans_36_leadingZeros_T_93[32] ? 6'h20 : _ans_36_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_159 = _ans_36_leadingZeros_T_93[31] ? 6'h1f : _ans_36_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_160 = _ans_36_leadingZeros_T_93[30] ? 6'h1e : _ans_36_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_161 = _ans_36_leadingZeros_T_93[29] ? 6'h1d : _ans_36_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_162 = _ans_36_leadingZeros_T_93[28] ? 6'h1c : _ans_36_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_163 = _ans_36_leadingZeros_T_93[27] ? 6'h1b : _ans_36_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_164 = _ans_36_leadingZeros_T_93[26] ? 6'h1a : _ans_36_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_165 = _ans_36_leadingZeros_T_93[25] ? 6'h19 : _ans_36_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_166 = _ans_36_leadingZeros_T_93[24] ? 6'h18 : _ans_36_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_167 = _ans_36_leadingZeros_T_93[23] ? 6'h17 : _ans_36_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_168 = _ans_36_leadingZeros_T_93[22] ? 6'h16 : _ans_36_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_169 = _ans_36_leadingZeros_T_93[21] ? 6'h15 : _ans_36_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_170 = _ans_36_leadingZeros_T_93[20] ? 6'h14 : _ans_36_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_171 = _ans_36_leadingZeros_T_93[19] ? 6'h13 : _ans_36_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_172 = _ans_36_leadingZeros_T_93[18] ? 6'h12 : _ans_36_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_173 = _ans_36_leadingZeros_T_93[17] ? 6'h11 : _ans_36_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_174 = _ans_36_leadingZeros_T_93[16] ? 6'h10 : _ans_36_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_175 = _ans_36_leadingZeros_T_93[15] ? 6'hf : _ans_36_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_176 = _ans_36_leadingZeros_T_93[14] ? 6'he : _ans_36_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_177 = _ans_36_leadingZeros_T_93[13] ? 6'hd : _ans_36_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_178 = _ans_36_leadingZeros_T_93[12] ? 6'hc : _ans_36_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_179 = _ans_36_leadingZeros_T_93[11] ? 6'hb : _ans_36_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_180 = _ans_36_leadingZeros_T_93[10] ? 6'ha : _ans_36_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_181 = _ans_36_leadingZeros_T_93[9] ? 6'h9 : _ans_36_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_182 = _ans_36_leadingZeros_T_93[8] ? 6'h8 : _ans_36_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_183 = _ans_36_leadingZeros_T_93[7] ? 6'h7 : _ans_36_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_184 = _ans_36_leadingZeros_T_93[6] ? 6'h6 : _ans_36_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_185 = _ans_36_leadingZeros_T_93[5] ? 6'h5 : _ans_36_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_186 = _ans_36_leadingZeros_T_93[4] ? 6'h4 : _ans_36_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_187 = _ans_36_leadingZeros_T_93[3] ? 6'h3 : _ans_36_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_188 = _ans_36_leadingZeros_T_93[2] ? 6'h2 : _ans_36_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_leadingZeros_T_189 = _ans_36_leadingZeros_T_93[1] ? 6'h1 : _ans_36_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_36_leadingZeros = _ans_36_leadingZeros_T_93[0] ? 6'h0 : _ans_36_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_36_expRaw_T_1 = 6'h1f - ans_36_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_36_expRaw = ans_36_isZero ? 6'h0 : _ans_36_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_36_shiftAmt_T_2 = ans_36_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_36_shiftAmt = ans_36_expRaw > 6'h3 ? _ans_36_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_36_mantissaRaw_T = ans_36_absClipped >> ans_36_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_36_mantissaRaw = _ans_36_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_36_mantissa = ans_36_expRaw >= 6'h3 ? ans_36_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_36_expAdjusted = ans_36_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_36_exp_T_4 = ans_36_expAdjusted > 7'hf ? 4'hf : ans_36_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_36_exp = ans_36_isZero ? 4'h0 : _ans_36_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_36_fp8 = {ans_36_clippedX[31],ans_36_exp,ans_36_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_37 = {24'h0,linear_bias_37}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_37 = tempSum_37 + biasExtended_37; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_37_sign = sum32_37[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_37_absX_T = ~sum32_37; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_37_absX_T_2 = _ans_37_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_37_absX = ans_37_sign ? _ans_37_absX_T_2 : sum32_37; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_37_shiftedX_T_1 = _GEN_10432 - ans_37_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_37_shiftedX_T_3 = ans_37_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_37_shiftedX = ans_37_sign ? _ans_37_shiftedX_T_1 : _ans_37_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_37_scaledX_T_1 = ans_37_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_37_scaledX = _ans_37_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_37_clippedX_T_2 = ans_37_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_37_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_37_clippedX = ans_37_scaledX > 49'h1c0 ? 49'h1c0 : _ans_37_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_37_absClipped_T_1 = ~ans_37_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_37_absClipped_T_3 = _ans_37_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_37_absClipped = ans_37_clippedX[31] ? _ans_37_absClipped_T_3 : ans_37_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_37_isZero = ans_37_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10841 = {{16'd0}, ans_37_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_4 = _GEN_10841 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_6 = {ans_37_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_8 = _ans_37_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_9 = _ans_37_leadingZeros_T_4 | _ans_37_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10842 = {{8'd0}, _ans_37_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_14 = _GEN_10842 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_16 = {_ans_37_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_18 = _ans_37_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_19 = _ans_37_leadingZeros_T_14 | _ans_37_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10843 = {{4'd0}, _ans_37_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_24 = _GEN_10843 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_26 = {_ans_37_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_28 = _ans_37_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_29 = _ans_37_leadingZeros_T_24 | _ans_37_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10844 = {{2'd0}, _ans_37_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_34 = _GEN_10844 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_36 = {_ans_37_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_38 = _ans_37_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_39 = _ans_37_leadingZeros_T_34 | _ans_37_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10845 = {{1'd0}, _ans_37_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_44 = _GEN_10845 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_46 = {_ans_37_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_48 = _ans_37_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_37_leadingZeros_T_49 = _ans_37_leadingZeros_T_44 | _ans_37_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10846 = {{8'd0}, ans_37_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_55 = _GEN_10846 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_57 = {ans_37_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_59 = _ans_37_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_60 = _ans_37_leadingZeros_T_55 | _ans_37_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10847 = {{4'd0}, _ans_37_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_65 = _GEN_10847 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_67 = {_ans_37_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_69 = _ans_37_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_70 = _ans_37_leadingZeros_T_65 | _ans_37_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10848 = {{2'd0}, _ans_37_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_75 = _GEN_10848 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_77 = {_ans_37_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_79 = _ans_37_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_80 = _ans_37_leadingZeros_T_75 | _ans_37_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10849 = {{1'd0}, _ans_37_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_85 = _GEN_10849 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_87 = {_ans_37_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_89 = _ans_37_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_37_leadingZeros_T_90 = _ans_37_leadingZeros_T_85 | _ans_37_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_37_leadingZeros_T_93 = {_ans_37_leadingZeros_T_49,_ans_37_leadingZeros_T_90,ans_37_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_37_leadingZeros_T_143 = _ans_37_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_144 = _ans_37_leadingZeros_T_93[46] ? 6'h2e : _ans_37_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_145 = _ans_37_leadingZeros_T_93[45] ? 6'h2d : _ans_37_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_146 = _ans_37_leadingZeros_T_93[44] ? 6'h2c : _ans_37_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_147 = _ans_37_leadingZeros_T_93[43] ? 6'h2b : _ans_37_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_148 = _ans_37_leadingZeros_T_93[42] ? 6'h2a : _ans_37_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_149 = _ans_37_leadingZeros_T_93[41] ? 6'h29 : _ans_37_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_150 = _ans_37_leadingZeros_T_93[40] ? 6'h28 : _ans_37_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_151 = _ans_37_leadingZeros_T_93[39] ? 6'h27 : _ans_37_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_152 = _ans_37_leadingZeros_T_93[38] ? 6'h26 : _ans_37_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_153 = _ans_37_leadingZeros_T_93[37] ? 6'h25 : _ans_37_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_154 = _ans_37_leadingZeros_T_93[36] ? 6'h24 : _ans_37_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_155 = _ans_37_leadingZeros_T_93[35] ? 6'h23 : _ans_37_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_156 = _ans_37_leadingZeros_T_93[34] ? 6'h22 : _ans_37_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_157 = _ans_37_leadingZeros_T_93[33] ? 6'h21 : _ans_37_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_158 = _ans_37_leadingZeros_T_93[32] ? 6'h20 : _ans_37_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_159 = _ans_37_leadingZeros_T_93[31] ? 6'h1f : _ans_37_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_160 = _ans_37_leadingZeros_T_93[30] ? 6'h1e : _ans_37_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_161 = _ans_37_leadingZeros_T_93[29] ? 6'h1d : _ans_37_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_162 = _ans_37_leadingZeros_T_93[28] ? 6'h1c : _ans_37_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_163 = _ans_37_leadingZeros_T_93[27] ? 6'h1b : _ans_37_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_164 = _ans_37_leadingZeros_T_93[26] ? 6'h1a : _ans_37_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_165 = _ans_37_leadingZeros_T_93[25] ? 6'h19 : _ans_37_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_166 = _ans_37_leadingZeros_T_93[24] ? 6'h18 : _ans_37_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_167 = _ans_37_leadingZeros_T_93[23] ? 6'h17 : _ans_37_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_168 = _ans_37_leadingZeros_T_93[22] ? 6'h16 : _ans_37_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_169 = _ans_37_leadingZeros_T_93[21] ? 6'h15 : _ans_37_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_170 = _ans_37_leadingZeros_T_93[20] ? 6'h14 : _ans_37_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_171 = _ans_37_leadingZeros_T_93[19] ? 6'h13 : _ans_37_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_172 = _ans_37_leadingZeros_T_93[18] ? 6'h12 : _ans_37_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_173 = _ans_37_leadingZeros_T_93[17] ? 6'h11 : _ans_37_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_174 = _ans_37_leadingZeros_T_93[16] ? 6'h10 : _ans_37_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_175 = _ans_37_leadingZeros_T_93[15] ? 6'hf : _ans_37_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_176 = _ans_37_leadingZeros_T_93[14] ? 6'he : _ans_37_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_177 = _ans_37_leadingZeros_T_93[13] ? 6'hd : _ans_37_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_178 = _ans_37_leadingZeros_T_93[12] ? 6'hc : _ans_37_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_179 = _ans_37_leadingZeros_T_93[11] ? 6'hb : _ans_37_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_180 = _ans_37_leadingZeros_T_93[10] ? 6'ha : _ans_37_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_181 = _ans_37_leadingZeros_T_93[9] ? 6'h9 : _ans_37_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_182 = _ans_37_leadingZeros_T_93[8] ? 6'h8 : _ans_37_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_183 = _ans_37_leadingZeros_T_93[7] ? 6'h7 : _ans_37_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_184 = _ans_37_leadingZeros_T_93[6] ? 6'h6 : _ans_37_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_185 = _ans_37_leadingZeros_T_93[5] ? 6'h5 : _ans_37_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_186 = _ans_37_leadingZeros_T_93[4] ? 6'h4 : _ans_37_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_187 = _ans_37_leadingZeros_T_93[3] ? 6'h3 : _ans_37_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_188 = _ans_37_leadingZeros_T_93[2] ? 6'h2 : _ans_37_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_leadingZeros_T_189 = _ans_37_leadingZeros_T_93[1] ? 6'h1 : _ans_37_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_37_leadingZeros = _ans_37_leadingZeros_T_93[0] ? 6'h0 : _ans_37_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_37_expRaw_T_1 = 6'h1f - ans_37_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_37_expRaw = ans_37_isZero ? 6'h0 : _ans_37_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_37_shiftAmt_T_2 = ans_37_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_37_shiftAmt = ans_37_expRaw > 6'h3 ? _ans_37_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_37_mantissaRaw_T = ans_37_absClipped >> ans_37_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_37_mantissaRaw = _ans_37_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_37_mantissa = ans_37_expRaw >= 6'h3 ? ans_37_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_37_expAdjusted = ans_37_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_37_exp_T_4 = ans_37_expAdjusted > 7'hf ? 4'hf : ans_37_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_37_exp = ans_37_isZero ? 4'h0 : _ans_37_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_37_fp8 = {ans_37_clippedX[31],ans_37_exp,ans_37_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_38 = {24'h0,linear_bias_38}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_38 = tempSum_38 + biasExtended_38; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_38_sign = sum32_38[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_38_absX_T = ~sum32_38; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_38_absX_T_2 = _ans_38_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_38_absX = ans_38_sign ? _ans_38_absX_T_2 : sum32_38; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_38_shiftedX_T_1 = _GEN_10432 - ans_38_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_38_shiftedX_T_3 = ans_38_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_38_shiftedX = ans_38_sign ? _ans_38_shiftedX_T_1 : _ans_38_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_38_scaledX_T_1 = ans_38_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_38_scaledX = _ans_38_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_38_clippedX_T_2 = ans_38_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_38_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_38_clippedX = ans_38_scaledX > 49'h1c0 ? 49'h1c0 : _ans_38_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_38_absClipped_T_1 = ~ans_38_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_38_absClipped_T_3 = _ans_38_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_38_absClipped = ans_38_clippedX[31] ? _ans_38_absClipped_T_3 : ans_38_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_38_isZero = ans_38_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10852 = {{16'd0}, ans_38_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_4 = _GEN_10852 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_6 = {ans_38_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_8 = _ans_38_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_9 = _ans_38_leadingZeros_T_4 | _ans_38_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10853 = {{8'd0}, _ans_38_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_14 = _GEN_10853 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_16 = {_ans_38_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_18 = _ans_38_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_19 = _ans_38_leadingZeros_T_14 | _ans_38_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10854 = {{4'd0}, _ans_38_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_24 = _GEN_10854 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_26 = {_ans_38_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_28 = _ans_38_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_29 = _ans_38_leadingZeros_T_24 | _ans_38_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10855 = {{2'd0}, _ans_38_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_34 = _GEN_10855 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_36 = {_ans_38_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_38 = _ans_38_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_39 = _ans_38_leadingZeros_T_34 | _ans_38_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10856 = {{1'd0}, _ans_38_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_44 = _GEN_10856 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_46 = {_ans_38_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_48 = _ans_38_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_38_leadingZeros_T_49 = _ans_38_leadingZeros_T_44 | _ans_38_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10857 = {{8'd0}, ans_38_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_55 = _GEN_10857 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_57 = {ans_38_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_59 = _ans_38_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_60 = _ans_38_leadingZeros_T_55 | _ans_38_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10858 = {{4'd0}, _ans_38_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_65 = _GEN_10858 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_67 = {_ans_38_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_69 = _ans_38_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_70 = _ans_38_leadingZeros_T_65 | _ans_38_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10859 = {{2'd0}, _ans_38_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_75 = _GEN_10859 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_77 = {_ans_38_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_79 = _ans_38_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_80 = _ans_38_leadingZeros_T_75 | _ans_38_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10860 = {{1'd0}, _ans_38_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_85 = _GEN_10860 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_87 = {_ans_38_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_89 = _ans_38_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_38_leadingZeros_T_90 = _ans_38_leadingZeros_T_85 | _ans_38_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_38_leadingZeros_T_93 = {_ans_38_leadingZeros_T_49,_ans_38_leadingZeros_T_90,ans_38_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_38_leadingZeros_T_143 = _ans_38_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_144 = _ans_38_leadingZeros_T_93[46] ? 6'h2e : _ans_38_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_145 = _ans_38_leadingZeros_T_93[45] ? 6'h2d : _ans_38_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_146 = _ans_38_leadingZeros_T_93[44] ? 6'h2c : _ans_38_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_147 = _ans_38_leadingZeros_T_93[43] ? 6'h2b : _ans_38_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_148 = _ans_38_leadingZeros_T_93[42] ? 6'h2a : _ans_38_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_149 = _ans_38_leadingZeros_T_93[41] ? 6'h29 : _ans_38_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_150 = _ans_38_leadingZeros_T_93[40] ? 6'h28 : _ans_38_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_151 = _ans_38_leadingZeros_T_93[39] ? 6'h27 : _ans_38_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_152 = _ans_38_leadingZeros_T_93[38] ? 6'h26 : _ans_38_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_153 = _ans_38_leadingZeros_T_93[37] ? 6'h25 : _ans_38_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_154 = _ans_38_leadingZeros_T_93[36] ? 6'h24 : _ans_38_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_155 = _ans_38_leadingZeros_T_93[35] ? 6'h23 : _ans_38_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_156 = _ans_38_leadingZeros_T_93[34] ? 6'h22 : _ans_38_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_157 = _ans_38_leadingZeros_T_93[33] ? 6'h21 : _ans_38_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_158 = _ans_38_leadingZeros_T_93[32] ? 6'h20 : _ans_38_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_159 = _ans_38_leadingZeros_T_93[31] ? 6'h1f : _ans_38_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_160 = _ans_38_leadingZeros_T_93[30] ? 6'h1e : _ans_38_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_161 = _ans_38_leadingZeros_T_93[29] ? 6'h1d : _ans_38_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_162 = _ans_38_leadingZeros_T_93[28] ? 6'h1c : _ans_38_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_163 = _ans_38_leadingZeros_T_93[27] ? 6'h1b : _ans_38_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_164 = _ans_38_leadingZeros_T_93[26] ? 6'h1a : _ans_38_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_165 = _ans_38_leadingZeros_T_93[25] ? 6'h19 : _ans_38_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_166 = _ans_38_leadingZeros_T_93[24] ? 6'h18 : _ans_38_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_167 = _ans_38_leadingZeros_T_93[23] ? 6'h17 : _ans_38_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_168 = _ans_38_leadingZeros_T_93[22] ? 6'h16 : _ans_38_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_169 = _ans_38_leadingZeros_T_93[21] ? 6'h15 : _ans_38_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_170 = _ans_38_leadingZeros_T_93[20] ? 6'h14 : _ans_38_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_171 = _ans_38_leadingZeros_T_93[19] ? 6'h13 : _ans_38_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_172 = _ans_38_leadingZeros_T_93[18] ? 6'h12 : _ans_38_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_173 = _ans_38_leadingZeros_T_93[17] ? 6'h11 : _ans_38_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_174 = _ans_38_leadingZeros_T_93[16] ? 6'h10 : _ans_38_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_175 = _ans_38_leadingZeros_T_93[15] ? 6'hf : _ans_38_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_176 = _ans_38_leadingZeros_T_93[14] ? 6'he : _ans_38_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_177 = _ans_38_leadingZeros_T_93[13] ? 6'hd : _ans_38_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_178 = _ans_38_leadingZeros_T_93[12] ? 6'hc : _ans_38_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_179 = _ans_38_leadingZeros_T_93[11] ? 6'hb : _ans_38_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_180 = _ans_38_leadingZeros_T_93[10] ? 6'ha : _ans_38_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_181 = _ans_38_leadingZeros_T_93[9] ? 6'h9 : _ans_38_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_182 = _ans_38_leadingZeros_T_93[8] ? 6'h8 : _ans_38_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_183 = _ans_38_leadingZeros_T_93[7] ? 6'h7 : _ans_38_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_184 = _ans_38_leadingZeros_T_93[6] ? 6'h6 : _ans_38_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_185 = _ans_38_leadingZeros_T_93[5] ? 6'h5 : _ans_38_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_186 = _ans_38_leadingZeros_T_93[4] ? 6'h4 : _ans_38_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_187 = _ans_38_leadingZeros_T_93[3] ? 6'h3 : _ans_38_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_188 = _ans_38_leadingZeros_T_93[2] ? 6'h2 : _ans_38_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_leadingZeros_T_189 = _ans_38_leadingZeros_T_93[1] ? 6'h1 : _ans_38_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_38_leadingZeros = _ans_38_leadingZeros_T_93[0] ? 6'h0 : _ans_38_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_38_expRaw_T_1 = 6'h1f - ans_38_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_38_expRaw = ans_38_isZero ? 6'h0 : _ans_38_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_38_shiftAmt_T_2 = ans_38_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_38_shiftAmt = ans_38_expRaw > 6'h3 ? _ans_38_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_38_mantissaRaw_T = ans_38_absClipped >> ans_38_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_38_mantissaRaw = _ans_38_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_38_mantissa = ans_38_expRaw >= 6'h3 ? ans_38_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_38_expAdjusted = ans_38_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_38_exp_T_4 = ans_38_expAdjusted > 7'hf ? 4'hf : ans_38_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_38_exp = ans_38_isZero ? 4'h0 : _ans_38_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_38_fp8 = {ans_38_clippedX[31],ans_38_exp,ans_38_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_39 = {24'h0,linear_bias_39}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_39 = tempSum_39 + biasExtended_39; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_39_sign = sum32_39[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_39_absX_T = ~sum32_39; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_39_absX_T_2 = _ans_39_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_39_absX = ans_39_sign ? _ans_39_absX_T_2 : sum32_39; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_39_shiftedX_T_1 = _GEN_10432 - ans_39_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_39_shiftedX_T_3 = ans_39_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_39_shiftedX = ans_39_sign ? _ans_39_shiftedX_T_1 : _ans_39_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_39_scaledX_T_1 = ans_39_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_39_scaledX = _ans_39_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_39_clippedX_T_2 = ans_39_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_39_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_39_clippedX = ans_39_scaledX > 49'h1c0 ? 49'h1c0 : _ans_39_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_39_absClipped_T_1 = ~ans_39_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_39_absClipped_T_3 = _ans_39_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_39_absClipped = ans_39_clippedX[31] ? _ans_39_absClipped_T_3 : ans_39_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_39_isZero = ans_39_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10863 = {{16'd0}, ans_39_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_4 = _GEN_10863 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_6 = {ans_39_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_8 = _ans_39_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_9 = _ans_39_leadingZeros_T_4 | _ans_39_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10864 = {{8'd0}, _ans_39_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_14 = _GEN_10864 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_16 = {_ans_39_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_18 = _ans_39_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_19 = _ans_39_leadingZeros_T_14 | _ans_39_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10865 = {{4'd0}, _ans_39_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_24 = _GEN_10865 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_26 = {_ans_39_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_28 = _ans_39_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_29 = _ans_39_leadingZeros_T_24 | _ans_39_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10866 = {{2'd0}, _ans_39_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_34 = _GEN_10866 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_36 = {_ans_39_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_38 = _ans_39_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_39 = _ans_39_leadingZeros_T_34 | _ans_39_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10867 = {{1'd0}, _ans_39_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_44 = _GEN_10867 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_46 = {_ans_39_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_48 = _ans_39_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_39_leadingZeros_T_49 = _ans_39_leadingZeros_T_44 | _ans_39_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10868 = {{8'd0}, ans_39_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_55 = _GEN_10868 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_57 = {ans_39_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_59 = _ans_39_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_60 = _ans_39_leadingZeros_T_55 | _ans_39_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10869 = {{4'd0}, _ans_39_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_65 = _GEN_10869 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_67 = {_ans_39_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_69 = _ans_39_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_70 = _ans_39_leadingZeros_T_65 | _ans_39_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10870 = {{2'd0}, _ans_39_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_75 = _GEN_10870 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_77 = {_ans_39_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_79 = _ans_39_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_80 = _ans_39_leadingZeros_T_75 | _ans_39_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10871 = {{1'd0}, _ans_39_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_85 = _GEN_10871 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_87 = {_ans_39_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_89 = _ans_39_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_39_leadingZeros_T_90 = _ans_39_leadingZeros_T_85 | _ans_39_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_39_leadingZeros_T_93 = {_ans_39_leadingZeros_T_49,_ans_39_leadingZeros_T_90,ans_39_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_39_leadingZeros_T_143 = _ans_39_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_144 = _ans_39_leadingZeros_T_93[46] ? 6'h2e : _ans_39_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_145 = _ans_39_leadingZeros_T_93[45] ? 6'h2d : _ans_39_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_146 = _ans_39_leadingZeros_T_93[44] ? 6'h2c : _ans_39_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_147 = _ans_39_leadingZeros_T_93[43] ? 6'h2b : _ans_39_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_148 = _ans_39_leadingZeros_T_93[42] ? 6'h2a : _ans_39_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_149 = _ans_39_leadingZeros_T_93[41] ? 6'h29 : _ans_39_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_150 = _ans_39_leadingZeros_T_93[40] ? 6'h28 : _ans_39_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_151 = _ans_39_leadingZeros_T_93[39] ? 6'h27 : _ans_39_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_152 = _ans_39_leadingZeros_T_93[38] ? 6'h26 : _ans_39_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_153 = _ans_39_leadingZeros_T_93[37] ? 6'h25 : _ans_39_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_154 = _ans_39_leadingZeros_T_93[36] ? 6'h24 : _ans_39_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_155 = _ans_39_leadingZeros_T_93[35] ? 6'h23 : _ans_39_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_156 = _ans_39_leadingZeros_T_93[34] ? 6'h22 : _ans_39_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_157 = _ans_39_leadingZeros_T_93[33] ? 6'h21 : _ans_39_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_158 = _ans_39_leadingZeros_T_93[32] ? 6'h20 : _ans_39_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_159 = _ans_39_leadingZeros_T_93[31] ? 6'h1f : _ans_39_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_160 = _ans_39_leadingZeros_T_93[30] ? 6'h1e : _ans_39_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_161 = _ans_39_leadingZeros_T_93[29] ? 6'h1d : _ans_39_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_162 = _ans_39_leadingZeros_T_93[28] ? 6'h1c : _ans_39_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_163 = _ans_39_leadingZeros_T_93[27] ? 6'h1b : _ans_39_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_164 = _ans_39_leadingZeros_T_93[26] ? 6'h1a : _ans_39_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_165 = _ans_39_leadingZeros_T_93[25] ? 6'h19 : _ans_39_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_166 = _ans_39_leadingZeros_T_93[24] ? 6'h18 : _ans_39_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_167 = _ans_39_leadingZeros_T_93[23] ? 6'h17 : _ans_39_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_168 = _ans_39_leadingZeros_T_93[22] ? 6'h16 : _ans_39_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_169 = _ans_39_leadingZeros_T_93[21] ? 6'h15 : _ans_39_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_170 = _ans_39_leadingZeros_T_93[20] ? 6'h14 : _ans_39_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_171 = _ans_39_leadingZeros_T_93[19] ? 6'h13 : _ans_39_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_172 = _ans_39_leadingZeros_T_93[18] ? 6'h12 : _ans_39_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_173 = _ans_39_leadingZeros_T_93[17] ? 6'h11 : _ans_39_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_174 = _ans_39_leadingZeros_T_93[16] ? 6'h10 : _ans_39_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_175 = _ans_39_leadingZeros_T_93[15] ? 6'hf : _ans_39_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_176 = _ans_39_leadingZeros_T_93[14] ? 6'he : _ans_39_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_177 = _ans_39_leadingZeros_T_93[13] ? 6'hd : _ans_39_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_178 = _ans_39_leadingZeros_T_93[12] ? 6'hc : _ans_39_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_179 = _ans_39_leadingZeros_T_93[11] ? 6'hb : _ans_39_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_180 = _ans_39_leadingZeros_T_93[10] ? 6'ha : _ans_39_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_181 = _ans_39_leadingZeros_T_93[9] ? 6'h9 : _ans_39_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_182 = _ans_39_leadingZeros_T_93[8] ? 6'h8 : _ans_39_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_183 = _ans_39_leadingZeros_T_93[7] ? 6'h7 : _ans_39_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_184 = _ans_39_leadingZeros_T_93[6] ? 6'h6 : _ans_39_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_185 = _ans_39_leadingZeros_T_93[5] ? 6'h5 : _ans_39_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_186 = _ans_39_leadingZeros_T_93[4] ? 6'h4 : _ans_39_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_187 = _ans_39_leadingZeros_T_93[3] ? 6'h3 : _ans_39_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_188 = _ans_39_leadingZeros_T_93[2] ? 6'h2 : _ans_39_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_leadingZeros_T_189 = _ans_39_leadingZeros_T_93[1] ? 6'h1 : _ans_39_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_39_leadingZeros = _ans_39_leadingZeros_T_93[0] ? 6'h0 : _ans_39_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_39_expRaw_T_1 = 6'h1f - ans_39_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_39_expRaw = ans_39_isZero ? 6'h0 : _ans_39_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_39_shiftAmt_T_2 = ans_39_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_39_shiftAmt = ans_39_expRaw > 6'h3 ? _ans_39_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_39_mantissaRaw_T = ans_39_absClipped >> ans_39_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_39_mantissaRaw = _ans_39_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_39_mantissa = ans_39_expRaw >= 6'h3 ? ans_39_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_39_expAdjusted = ans_39_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_39_exp_T_4 = ans_39_expAdjusted > 7'hf ? 4'hf : ans_39_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_39_exp = ans_39_isZero ? 4'h0 : _ans_39_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_39_fp8 = {ans_39_clippedX[31],ans_39_exp,ans_39_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_40 = {24'h0,linear_bias_40}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_40 = tempSum_40 + biasExtended_40; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_40_sign = sum32_40[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_40_absX_T = ~sum32_40; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_40_absX_T_2 = _ans_40_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_40_absX = ans_40_sign ? _ans_40_absX_T_2 : sum32_40; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_40_shiftedX_T_1 = _GEN_10432 - ans_40_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_40_shiftedX_T_3 = ans_40_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_40_shiftedX = ans_40_sign ? _ans_40_shiftedX_T_1 : _ans_40_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_40_scaledX_T_1 = ans_40_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_40_scaledX = _ans_40_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_40_clippedX_T_2 = ans_40_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_40_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_40_clippedX = ans_40_scaledX > 49'h1c0 ? 49'h1c0 : _ans_40_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_40_absClipped_T_1 = ~ans_40_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_40_absClipped_T_3 = _ans_40_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_40_absClipped = ans_40_clippedX[31] ? _ans_40_absClipped_T_3 : ans_40_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_40_isZero = ans_40_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10874 = {{16'd0}, ans_40_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_4 = _GEN_10874 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_6 = {ans_40_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_8 = _ans_40_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_9 = _ans_40_leadingZeros_T_4 | _ans_40_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10875 = {{8'd0}, _ans_40_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_14 = _GEN_10875 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_16 = {_ans_40_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_18 = _ans_40_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_19 = _ans_40_leadingZeros_T_14 | _ans_40_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10876 = {{4'd0}, _ans_40_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_24 = _GEN_10876 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_26 = {_ans_40_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_28 = _ans_40_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_29 = _ans_40_leadingZeros_T_24 | _ans_40_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10877 = {{2'd0}, _ans_40_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_34 = _GEN_10877 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_36 = {_ans_40_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_38 = _ans_40_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_39 = _ans_40_leadingZeros_T_34 | _ans_40_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10878 = {{1'd0}, _ans_40_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_44 = _GEN_10878 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_46 = {_ans_40_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_48 = _ans_40_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_40_leadingZeros_T_49 = _ans_40_leadingZeros_T_44 | _ans_40_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10879 = {{8'd0}, ans_40_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_55 = _GEN_10879 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_57 = {ans_40_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_59 = _ans_40_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_60 = _ans_40_leadingZeros_T_55 | _ans_40_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10880 = {{4'd0}, _ans_40_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_65 = _GEN_10880 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_67 = {_ans_40_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_69 = _ans_40_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_70 = _ans_40_leadingZeros_T_65 | _ans_40_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10881 = {{2'd0}, _ans_40_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_75 = _GEN_10881 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_77 = {_ans_40_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_79 = _ans_40_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_80 = _ans_40_leadingZeros_T_75 | _ans_40_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10882 = {{1'd0}, _ans_40_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_85 = _GEN_10882 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_87 = {_ans_40_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_89 = _ans_40_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_40_leadingZeros_T_90 = _ans_40_leadingZeros_T_85 | _ans_40_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_40_leadingZeros_T_93 = {_ans_40_leadingZeros_T_49,_ans_40_leadingZeros_T_90,ans_40_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_40_leadingZeros_T_143 = _ans_40_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_144 = _ans_40_leadingZeros_T_93[46] ? 6'h2e : _ans_40_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_145 = _ans_40_leadingZeros_T_93[45] ? 6'h2d : _ans_40_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_146 = _ans_40_leadingZeros_T_93[44] ? 6'h2c : _ans_40_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_147 = _ans_40_leadingZeros_T_93[43] ? 6'h2b : _ans_40_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_148 = _ans_40_leadingZeros_T_93[42] ? 6'h2a : _ans_40_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_149 = _ans_40_leadingZeros_T_93[41] ? 6'h29 : _ans_40_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_150 = _ans_40_leadingZeros_T_93[40] ? 6'h28 : _ans_40_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_151 = _ans_40_leadingZeros_T_93[39] ? 6'h27 : _ans_40_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_152 = _ans_40_leadingZeros_T_93[38] ? 6'h26 : _ans_40_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_153 = _ans_40_leadingZeros_T_93[37] ? 6'h25 : _ans_40_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_154 = _ans_40_leadingZeros_T_93[36] ? 6'h24 : _ans_40_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_155 = _ans_40_leadingZeros_T_93[35] ? 6'h23 : _ans_40_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_156 = _ans_40_leadingZeros_T_93[34] ? 6'h22 : _ans_40_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_157 = _ans_40_leadingZeros_T_93[33] ? 6'h21 : _ans_40_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_158 = _ans_40_leadingZeros_T_93[32] ? 6'h20 : _ans_40_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_159 = _ans_40_leadingZeros_T_93[31] ? 6'h1f : _ans_40_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_160 = _ans_40_leadingZeros_T_93[30] ? 6'h1e : _ans_40_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_161 = _ans_40_leadingZeros_T_93[29] ? 6'h1d : _ans_40_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_162 = _ans_40_leadingZeros_T_93[28] ? 6'h1c : _ans_40_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_163 = _ans_40_leadingZeros_T_93[27] ? 6'h1b : _ans_40_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_164 = _ans_40_leadingZeros_T_93[26] ? 6'h1a : _ans_40_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_165 = _ans_40_leadingZeros_T_93[25] ? 6'h19 : _ans_40_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_166 = _ans_40_leadingZeros_T_93[24] ? 6'h18 : _ans_40_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_167 = _ans_40_leadingZeros_T_93[23] ? 6'h17 : _ans_40_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_168 = _ans_40_leadingZeros_T_93[22] ? 6'h16 : _ans_40_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_169 = _ans_40_leadingZeros_T_93[21] ? 6'h15 : _ans_40_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_170 = _ans_40_leadingZeros_T_93[20] ? 6'h14 : _ans_40_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_171 = _ans_40_leadingZeros_T_93[19] ? 6'h13 : _ans_40_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_172 = _ans_40_leadingZeros_T_93[18] ? 6'h12 : _ans_40_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_173 = _ans_40_leadingZeros_T_93[17] ? 6'h11 : _ans_40_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_174 = _ans_40_leadingZeros_T_93[16] ? 6'h10 : _ans_40_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_175 = _ans_40_leadingZeros_T_93[15] ? 6'hf : _ans_40_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_176 = _ans_40_leadingZeros_T_93[14] ? 6'he : _ans_40_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_177 = _ans_40_leadingZeros_T_93[13] ? 6'hd : _ans_40_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_178 = _ans_40_leadingZeros_T_93[12] ? 6'hc : _ans_40_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_179 = _ans_40_leadingZeros_T_93[11] ? 6'hb : _ans_40_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_180 = _ans_40_leadingZeros_T_93[10] ? 6'ha : _ans_40_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_181 = _ans_40_leadingZeros_T_93[9] ? 6'h9 : _ans_40_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_182 = _ans_40_leadingZeros_T_93[8] ? 6'h8 : _ans_40_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_183 = _ans_40_leadingZeros_T_93[7] ? 6'h7 : _ans_40_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_184 = _ans_40_leadingZeros_T_93[6] ? 6'h6 : _ans_40_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_185 = _ans_40_leadingZeros_T_93[5] ? 6'h5 : _ans_40_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_186 = _ans_40_leadingZeros_T_93[4] ? 6'h4 : _ans_40_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_187 = _ans_40_leadingZeros_T_93[3] ? 6'h3 : _ans_40_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_188 = _ans_40_leadingZeros_T_93[2] ? 6'h2 : _ans_40_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_leadingZeros_T_189 = _ans_40_leadingZeros_T_93[1] ? 6'h1 : _ans_40_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_40_leadingZeros = _ans_40_leadingZeros_T_93[0] ? 6'h0 : _ans_40_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_40_expRaw_T_1 = 6'h1f - ans_40_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_40_expRaw = ans_40_isZero ? 6'h0 : _ans_40_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_40_shiftAmt_T_2 = ans_40_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_40_shiftAmt = ans_40_expRaw > 6'h3 ? _ans_40_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_40_mantissaRaw_T = ans_40_absClipped >> ans_40_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_40_mantissaRaw = _ans_40_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_40_mantissa = ans_40_expRaw >= 6'h3 ? ans_40_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_40_expAdjusted = ans_40_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_40_exp_T_4 = ans_40_expAdjusted > 7'hf ? 4'hf : ans_40_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_40_exp = ans_40_isZero ? 4'h0 : _ans_40_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_40_fp8 = {ans_40_clippedX[31],ans_40_exp,ans_40_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_41 = {24'h0,linear_bias_41}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_41 = tempSum_41 + biasExtended_41; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_41_sign = sum32_41[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_41_absX_T = ~sum32_41; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_41_absX_T_2 = _ans_41_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_41_absX = ans_41_sign ? _ans_41_absX_T_2 : sum32_41; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_41_shiftedX_T_1 = _GEN_10432 - ans_41_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_41_shiftedX_T_3 = ans_41_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_41_shiftedX = ans_41_sign ? _ans_41_shiftedX_T_1 : _ans_41_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_41_scaledX_T_1 = ans_41_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_41_scaledX = _ans_41_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_41_clippedX_T_2 = ans_41_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_41_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_41_clippedX = ans_41_scaledX > 49'h1c0 ? 49'h1c0 : _ans_41_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_41_absClipped_T_1 = ~ans_41_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_41_absClipped_T_3 = _ans_41_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_41_absClipped = ans_41_clippedX[31] ? _ans_41_absClipped_T_3 : ans_41_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_41_isZero = ans_41_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10885 = {{16'd0}, ans_41_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_4 = _GEN_10885 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_6 = {ans_41_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_8 = _ans_41_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_9 = _ans_41_leadingZeros_T_4 | _ans_41_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10886 = {{8'd0}, _ans_41_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_14 = _GEN_10886 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_16 = {_ans_41_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_18 = _ans_41_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_19 = _ans_41_leadingZeros_T_14 | _ans_41_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10887 = {{4'd0}, _ans_41_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_24 = _GEN_10887 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_26 = {_ans_41_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_28 = _ans_41_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_29 = _ans_41_leadingZeros_T_24 | _ans_41_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10888 = {{2'd0}, _ans_41_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_34 = _GEN_10888 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_36 = {_ans_41_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_38 = _ans_41_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_39 = _ans_41_leadingZeros_T_34 | _ans_41_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10889 = {{1'd0}, _ans_41_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_44 = _GEN_10889 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_46 = {_ans_41_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_48 = _ans_41_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_41_leadingZeros_T_49 = _ans_41_leadingZeros_T_44 | _ans_41_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10890 = {{8'd0}, ans_41_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_55 = _GEN_10890 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_57 = {ans_41_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_59 = _ans_41_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_60 = _ans_41_leadingZeros_T_55 | _ans_41_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10891 = {{4'd0}, _ans_41_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_65 = _GEN_10891 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_67 = {_ans_41_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_69 = _ans_41_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_70 = _ans_41_leadingZeros_T_65 | _ans_41_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10892 = {{2'd0}, _ans_41_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_75 = _GEN_10892 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_77 = {_ans_41_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_79 = _ans_41_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_80 = _ans_41_leadingZeros_T_75 | _ans_41_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10893 = {{1'd0}, _ans_41_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_85 = _GEN_10893 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_87 = {_ans_41_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_89 = _ans_41_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_41_leadingZeros_T_90 = _ans_41_leadingZeros_T_85 | _ans_41_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_41_leadingZeros_T_93 = {_ans_41_leadingZeros_T_49,_ans_41_leadingZeros_T_90,ans_41_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_41_leadingZeros_T_143 = _ans_41_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_144 = _ans_41_leadingZeros_T_93[46] ? 6'h2e : _ans_41_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_145 = _ans_41_leadingZeros_T_93[45] ? 6'h2d : _ans_41_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_146 = _ans_41_leadingZeros_T_93[44] ? 6'h2c : _ans_41_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_147 = _ans_41_leadingZeros_T_93[43] ? 6'h2b : _ans_41_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_148 = _ans_41_leadingZeros_T_93[42] ? 6'h2a : _ans_41_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_149 = _ans_41_leadingZeros_T_93[41] ? 6'h29 : _ans_41_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_150 = _ans_41_leadingZeros_T_93[40] ? 6'h28 : _ans_41_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_151 = _ans_41_leadingZeros_T_93[39] ? 6'h27 : _ans_41_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_152 = _ans_41_leadingZeros_T_93[38] ? 6'h26 : _ans_41_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_153 = _ans_41_leadingZeros_T_93[37] ? 6'h25 : _ans_41_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_154 = _ans_41_leadingZeros_T_93[36] ? 6'h24 : _ans_41_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_155 = _ans_41_leadingZeros_T_93[35] ? 6'h23 : _ans_41_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_156 = _ans_41_leadingZeros_T_93[34] ? 6'h22 : _ans_41_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_157 = _ans_41_leadingZeros_T_93[33] ? 6'h21 : _ans_41_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_158 = _ans_41_leadingZeros_T_93[32] ? 6'h20 : _ans_41_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_159 = _ans_41_leadingZeros_T_93[31] ? 6'h1f : _ans_41_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_160 = _ans_41_leadingZeros_T_93[30] ? 6'h1e : _ans_41_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_161 = _ans_41_leadingZeros_T_93[29] ? 6'h1d : _ans_41_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_162 = _ans_41_leadingZeros_T_93[28] ? 6'h1c : _ans_41_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_163 = _ans_41_leadingZeros_T_93[27] ? 6'h1b : _ans_41_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_164 = _ans_41_leadingZeros_T_93[26] ? 6'h1a : _ans_41_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_165 = _ans_41_leadingZeros_T_93[25] ? 6'h19 : _ans_41_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_166 = _ans_41_leadingZeros_T_93[24] ? 6'h18 : _ans_41_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_167 = _ans_41_leadingZeros_T_93[23] ? 6'h17 : _ans_41_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_168 = _ans_41_leadingZeros_T_93[22] ? 6'h16 : _ans_41_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_169 = _ans_41_leadingZeros_T_93[21] ? 6'h15 : _ans_41_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_170 = _ans_41_leadingZeros_T_93[20] ? 6'h14 : _ans_41_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_171 = _ans_41_leadingZeros_T_93[19] ? 6'h13 : _ans_41_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_172 = _ans_41_leadingZeros_T_93[18] ? 6'h12 : _ans_41_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_173 = _ans_41_leadingZeros_T_93[17] ? 6'h11 : _ans_41_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_174 = _ans_41_leadingZeros_T_93[16] ? 6'h10 : _ans_41_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_175 = _ans_41_leadingZeros_T_93[15] ? 6'hf : _ans_41_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_176 = _ans_41_leadingZeros_T_93[14] ? 6'he : _ans_41_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_177 = _ans_41_leadingZeros_T_93[13] ? 6'hd : _ans_41_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_178 = _ans_41_leadingZeros_T_93[12] ? 6'hc : _ans_41_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_179 = _ans_41_leadingZeros_T_93[11] ? 6'hb : _ans_41_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_180 = _ans_41_leadingZeros_T_93[10] ? 6'ha : _ans_41_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_181 = _ans_41_leadingZeros_T_93[9] ? 6'h9 : _ans_41_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_182 = _ans_41_leadingZeros_T_93[8] ? 6'h8 : _ans_41_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_183 = _ans_41_leadingZeros_T_93[7] ? 6'h7 : _ans_41_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_184 = _ans_41_leadingZeros_T_93[6] ? 6'h6 : _ans_41_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_185 = _ans_41_leadingZeros_T_93[5] ? 6'h5 : _ans_41_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_186 = _ans_41_leadingZeros_T_93[4] ? 6'h4 : _ans_41_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_187 = _ans_41_leadingZeros_T_93[3] ? 6'h3 : _ans_41_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_188 = _ans_41_leadingZeros_T_93[2] ? 6'h2 : _ans_41_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_leadingZeros_T_189 = _ans_41_leadingZeros_T_93[1] ? 6'h1 : _ans_41_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_41_leadingZeros = _ans_41_leadingZeros_T_93[0] ? 6'h0 : _ans_41_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_41_expRaw_T_1 = 6'h1f - ans_41_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_41_expRaw = ans_41_isZero ? 6'h0 : _ans_41_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_41_shiftAmt_T_2 = ans_41_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_41_shiftAmt = ans_41_expRaw > 6'h3 ? _ans_41_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_41_mantissaRaw_T = ans_41_absClipped >> ans_41_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_41_mantissaRaw = _ans_41_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_41_mantissa = ans_41_expRaw >= 6'h3 ? ans_41_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_41_expAdjusted = ans_41_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_41_exp_T_4 = ans_41_expAdjusted > 7'hf ? 4'hf : ans_41_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_41_exp = ans_41_isZero ? 4'h0 : _ans_41_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_41_fp8 = {ans_41_clippedX[31],ans_41_exp,ans_41_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_42 = {24'h0,linear_bias_42}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_42 = tempSum_42 + biasExtended_42; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_42_sign = sum32_42[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_42_absX_T = ~sum32_42; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_42_absX_T_2 = _ans_42_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_42_absX = ans_42_sign ? _ans_42_absX_T_2 : sum32_42; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_42_shiftedX_T_1 = _GEN_10432 - ans_42_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_42_shiftedX_T_3 = ans_42_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_42_shiftedX = ans_42_sign ? _ans_42_shiftedX_T_1 : _ans_42_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_42_scaledX_T_1 = ans_42_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_42_scaledX = _ans_42_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_42_clippedX_T_2 = ans_42_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_42_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_42_clippedX = ans_42_scaledX > 49'h1c0 ? 49'h1c0 : _ans_42_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_42_absClipped_T_1 = ~ans_42_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_42_absClipped_T_3 = _ans_42_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_42_absClipped = ans_42_clippedX[31] ? _ans_42_absClipped_T_3 : ans_42_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_42_isZero = ans_42_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10896 = {{16'd0}, ans_42_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_4 = _GEN_10896 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_6 = {ans_42_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_8 = _ans_42_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_9 = _ans_42_leadingZeros_T_4 | _ans_42_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10897 = {{8'd0}, _ans_42_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_14 = _GEN_10897 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_16 = {_ans_42_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_18 = _ans_42_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_19 = _ans_42_leadingZeros_T_14 | _ans_42_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10898 = {{4'd0}, _ans_42_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_24 = _GEN_10898 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_26 = {_ans_42_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_28 = _ans_42_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_29 = _ans_42_leadingZeros_T_24 | _ans_42_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10899 = {{2'd0}, _ans_42_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_34 = _GEN_10899 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_36 = {_ans_42_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_38 = _ans_42_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_39 = _ans_42_leadingZeros_T_34 | _ans_42_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10900 = {{1'd0}, _ans_42_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_44 = _GEN_10900 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_46 = {_ans_42_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_48 = _ans_42_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_42_leadingZeros_T_49 = _ans_42_leadingZeros_T_44 | _ans_42_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10901 = {{8'd0}, ans_42_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_55 = _GEN_10901 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_57 = {ans_42_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_59 = _ans_42_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_60 = _ans_42_leadingZeros_T_55 | _ans_42_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10902 = {{4'd0}, _ans_42_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_65 = _GEN_10902 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_67 = {_ans_42_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_69 = _ans_42_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_70 = _ans_42_leadingZeros_T_65 | _ans_42_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10903 = {{2'd0}, _ans_42_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_75 = _GEN_10903 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_77 = {_ans_42_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_79 = _ans_42_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_80 = _ans_42_leadingZeros_T_75 | _ans_42_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10904 = {{1'd0}, _ans_42_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_85 = _GEN_10904 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_87 = {_ans_42_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_89 = _ans_42_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_42_leadingZeros_T_90 = _ans_42_leadingZeros_T_85 | _ans_42_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_42_leadingZeros_T_93 = {_ans_42_leadingZeros_T_49,_ans_42_leadingZeros_T_90,ans_42_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_42_leadingZeros_T_143 = _ans_42_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_144 = _ans_42_leadingZeros_T_93[46] ? 6'h2e : _ans_42_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_145 = _ans_42_leadingZeros_T_93[45] ? 6'h2d : _ans_42_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_146 = _ans_42_leadingZeros_T_93[44] ? 6'h2c : _ans_42_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_147 = _ans_42_leadingZeros_T_93[43] ? 6'h2b : _ans_42_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_148 = _ans_42_leadingZeros_T_93[42] ? 6'h2a : _ans_42_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_149 = _ans_42_leadingZeros_T_93[41] ? 6'h29 : _ans_42_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_150 = _ans_42_leadingZeros_T_93[40] ? 6'h28 : _ans_42_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_151 = _ans_42_leadingZeros_T_93[39] ? 6'h27 : _ans_42_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_152 = _ans_42_leadingZeros_T_93[38] ? 6'h26 : _ans_42_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_153 = _ans_42_leadingZeros_T_93[37] ? 6'h25 : _ans_42_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_154 = _ans_42_leadingZeros_T_93[36] ? 6'h24 : _ans_42_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_155 = _ans_42_leadingZeros_T_93[35] ? 6'h23 : _ans_42_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_156 = _ans_42_leadingZeros_T_93[34] ? 6'h22 : _ans_42_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_157 = _ans_42_leadingZeros_T_93[33] ? 6'h21 : _ans_42_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_158 = _ans_42_leadingZeros_T_93[32] ? 6'h20 : _ans_42_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_159 = _ans_42_leadingZeros_T_93[31] ? 6'h1f : _ans_42_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_160 = _ans_42_leadingZeros_T_93[30] ? 6'h1e : _ans_42_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_161 = _ans_42_leadingZeros_T_93[29] ? 6'h1d : _ans_42_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_162 = _ans_42_leadingZeros_T_93[28] ? 6'h1c : _ans_42_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_163 = _ans_42_leadingZeros_T_93[27] ? 6'h1b : _ans_42_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_164 = _ans_42_leadingZeros_T_93[26] ? 6'h1a : _ans_42_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_165 = _ans_42_leadingZeros_T_93[25] ? 6'h19 : _ans_42_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_166 = _ans_42_leadingZeros_T_93[24] ? 6'h18 : _ans_42_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_167 = _ans_42_leadingZeros_T_93[23] ? 6'h17 : _ans_42_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_168 = _ans_42_leadingZeros_T_93[22] ? 6'h16 : _ans_42_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_169 = _ans_42_leadingZeros_T_93[21] ? 6'h15 : _ans_42_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_170 = _ans_42_leadingZeros_T_93[20] ? 6'h14 : _ans_42_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_171 = _ans_42_leadingZeros_T_93[19] ? 6'h13 : _ans_42_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_172 = _ans_42_leadingZeros_T_93[18] ? 6'h12 : _ans_42_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_173 = _ans_42_leadingZeros_T_93[17] ? 6'h11 : _ans_42_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_174 = _ans_42_leadingZeros_T_93[16] ? 6'h10 : _ans_42_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_175 = _ans_42_leadingZeros_T_93[15] ? 6'hf : _ans_42_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_176 = _ans_42_leadingZeros_T_93[14] ? 6'he : _ans_42_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_177 = _ans_42_leadingZeros_T_93[13] ? 6'hd : _ans_42_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_178 = _ans_42_leadingZeros_T_93[12] ? 6'hc : _ans_42_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_179 = _ans_42_leadingZeros_T_93[11] ? 6'hb : _ans_42_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_180 = _ans_42_leadingZeros_T_93[10] ? 6'ha : _ans_42_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_181 = _ans_42_leadingZeros_T_93[9] ? 6'h9 : _ans_42_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_182 = _ans_42_leadingZeros_T_93[8] ? 6'h8 : _ans_42_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_183 = _ans_42_leadingZeros_T_93[7] ? 6'h7 : _ans_42_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_184 = _ans_42_leadingZeros_T_93[6] ? 6'h6 : _ans_42_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_185 = _ans_42_leadingZeros_T_93[5] ? 6'h5 : _ans_42_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_186 = _ans_42_leadingZeros_T_93[4] ? 6'h4 : _ans_42_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_187 = _ans_42_leadingZeros_T_93[3] ? 6'h3 : _ans_42_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_188 = _ans_42_leadingZeros_T_93[2] ? 6'h2 : _ans_42_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_leadingZeros_T_189 = _ans_42_leadingZeros_T_93[1] ? 6'h1 : _ans_42_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_42_leadingZeros = _ans_42_leadingZeros_T_93[0] ? 6'h0 : _ans_42_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_42_expRaw_T_1 = 6'h1f - ans_42_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_42_expRaw = ans_42_isZero ? 6'h0 : _ans_42_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_42_shiftAmt_T_2 = ans_42_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_42_shiftAmt = ans_42_expRaw > 6'h3 ? _ans_42_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_42_mantissaRaw_T = ans_42_absClipped >> ans_42_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_42_mantissaRaw = _ans_42_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_42_mantissa = ans_42_expRaw >= 6'h3 ? ans_42_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_42_expAdjusted = ans_42_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_42_exp_T_4 = ans_42_expAdjusted > 7'hf ? 4'hf : ans_42_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_42_exp = ans_42_isZero ? 4'h0 : _ans_42_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_42_fp8 = {ans_42_clippedX[31],ans_42_exp,ans_42_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_43 = {24'h0,linear_bias_43}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_43 = tempSum_43 + biasExtended_43; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_43_sign = sum32_43[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_43_absX_T = ~sum32_43; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_43_absX_T_2 = _ans_43_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_43_absX = ans_43_sign ? _ans_43_absX_T_2 : sum32_43; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_43_shiftedX_T_1 = _GEN_10432 - ans_43_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_43_shiftedX_T_3 = ans_43_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_43_shiftedX = ans_43_sign ? _ans_43_shiftedX_T_1 : _ans_43_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_43_scaledX_T_1 = ans_43_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_43_scaledX = _ans_43_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_43_clippedX_T_2 = ans_43_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_43_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_43_clippedX = ans_43_scaledX > 49'h1c0 ? 49'h1c0 : _ans_43_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_43_absClipped_T_1 = ~ans_43_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_43_absClipped_T_3 = _ans_43_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_43_absClipped = ans_43_clippedX[31] ? _ans_43_absClipped_T_3 : ans_43_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_43_isZero = ans_43_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10907 = {{16'd0}, ans_43_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_4 = _GEN_10907 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_6 = {ans_43_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_8 = _ans_43_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_9 = _ans_43_leadingZeros_T_4 | _ans_43_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10908 = {{8'd0}, _ans_43_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_14 = _GEN_10908 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_16 = {_ans_43_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_18 = _ans_43_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_19 = _ans_43_leadingZeros_T_14 | _ans_43_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10909 = {{4'd0}, _ans_43_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_24 = _GEN_10909 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_26 = {_ans_43_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_28 = _ans_43_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_29 = _ans_43_leadingZeros_T_24 | _ans_43_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10910 = {{2'd0}, _ans_43_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_34 = _GEN_10910 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_36 = {_ans_43_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_38 = _ans_43_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_39 = _ans_43_leadingZeros_T_34 | _ans_43_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10911 = {{1'd0}, _ans_43_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_44 = _GEN_10911 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_46 = {_ans_43_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_48 = _ans_43_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_43_leadingZeros_T_49 = _ans_43_leadingZeros_T_44 | _ans_43_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10912 = {{8'd0}, ans_43_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_55 = _GEN_10912 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_57 = {ans_43_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_59 = _ans_43_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_60 = _ans_43_leadingZeros_T_55 | _ans_43_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10913 = {{4'd0}, _ans_43_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_65 = _GEN_10913 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_67 = {_ans_43_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_69 = _ans_43_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_70 = _ans_43_leadingZeros_T_65 | _ans_43_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10914 = {{2'd0}, _ans_43_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_75 = _GEN_10914 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_77 = {_ans_43_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_79 = _ans_43_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_80 = _ans_43_leadingZeros_T_75 | _ans_43_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10915 = {{1'd0}, _ans_43_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_85 = _GEN_10915 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_87 = {_ans_43_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_89 = _ans_43_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_43_leadingZeros_T_90 = _ans_43_leadingZeros_T_85 | _ans_43_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_43_leadingZeros_T_93 = {_ans_43_leadingZeros_T_49,_ans_43_leadingZeros_T_90,ans_43_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_43_leadingZeros_T_143 = _ans_43_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_144 = _ans_43_leadingZeros_T_93[46] ? 6'h2e : _ans_43_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_145 = _ans_43_leadingZeros_T_93[45] ? 6'h2d : _ans_43_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_146 = _ans_43_leadingZeros_T_93[44] ? 6'h2c : _ans_43_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_147 = _ans_43_leadingZeros_T_93[43] ? 6'h2b : _ans_43_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_148 = _ans_43_leadingZeros_T_93[42] ? 6'h2a : _ans_43_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_149 = _ans_43_leadingZeros_T_93[41] ? 6'h29 : _ans_43_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_150 = _ans_43_leadingZeros_T_93[40] ? 6'h28 : _ans_43_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_151 = _ans_43_leadingZeros_T_93[39] ? 6'h27 : _ans_43_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_152 = _ans_43_leadingZeros_T_93[38] ? 6'h26 : _ans_43_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_153 = _ans_43_leadingZeros_T_93[37] ? 6'h25 : _ans_43_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_154 = _ans_43_leadingZeros_T_93[36] ? 6'h24 : _ans_43_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_155 = _ans_43_leadingZeros_T_93[35] ? 6'h23 : _ans_43_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_156 = _ans_43_leadingZeros_T_93[34] ? 6'h22 : _ans_43_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_157 = _ans_43_leadingZeros_T_93[33] ? 6'h21 : _ans_43_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_158 = _ans_43_leadingZeros_T_93[32] ? 6'h20 : _ans_43_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_159 = _ans_43_leadingZeros_T_93[31] ? 6'h1f : _ans_43_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_160 = _ans_43_leadingZeros_T_93[30] ? 6'h1e : _ans_43_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_161 = _ans_43_leadingZeros_T_93[29] ? 6'h1d : _ans_43_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_162 = _ans_43_leadingZeros_T_93[28] ? 6'h1c : _ans_43_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_163 = _ans_43_leadingZeros_T_93[27] ? 6'h1b : _ans_43_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_164 = _ans_43_leadingZeros_T_93[26] ? 6'h1a : _ans_43_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_165 = _ans_43_leadingZeros_T_93[25] ? 6'h19 : _ans_43_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_166 = _ans_43_leadingZeros_T_93[24] ? 6'h18 : _ans_43_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_167 = _ans_43_leadingZeros_T_93[23] ? 6'h17 : _ans_43_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_168 = _ans_43_leadingZeros_T_93[22] ? 6'h16 : _ans_43_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_169 = _ans_43_leadingZeros_T_93[21] ? 6'h15 : _ans_43_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_170 = _ans_43_leadingZeros_T_93[20] ? 6'h14 : _ans_43_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_171 = _ans_43_leadingZeros_T_93[19] ? 6'h13 : _ans_43_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_172 = _ans_43_leadingZeros_T_93[18] ? 6'h12 : _ans_43_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_173 = _ans_43_leadingZeros_T_93[17] ? 6'h11 : _ans_43_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_174 = _ans_43_leadingZeros_T_93[16] ? 6'h10 : _ans_43_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_175 = _ans_43_leadingZeros_T_93[15] ? 6'hf : _ans_43_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_176 = _ans_43_leadingZeros_T_93[14] ? 6'he : _ans_43_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_177 = _ans_43_leadingZeros_T_93[13] ? 6'hd : _ans_43_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_178 = _ans_43_leadingZeros_T_93[12] ? 6'hc : _ans_43_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_179 = _ans_43_leadingZeros_T_93[11] ? 6'hb : _ans_43_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_180 = _ans_43_leadingZeros_T_93[10] ? 6'ha : _ans_43_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_181 = _ans_43_leadingZeros_T_93[9] ? 6'h9 : _ans_43_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_182 = _ans_43_leadingZeros_T_93[8] ? 6'h8 : _ans_43_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_183 = _ans_43_leadingZeros_T_93[7] ? 6'h7 : _ans_43_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_184 = _ans_43_leadingZeros_T_93[6] ? 6'h6 : _ans_43_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_185 = _ans_43_leadingZeros_T_93[5] ? 6'h5 : _ans_43_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_186 = _ans_43_leadingZeros_T_93[4] ? 6'h4 : _ans_43_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_187 = _ans_43_leadingZeros_T_93[3] ? 6'h3 : _ans_43_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_188 = _ans_43_leadingZeros_T_93[2] ? 6'h2 : _ans_43_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_leadingZeros_T_189 = _ans_43_leadingZeros_T_93[1] ? 6'h1 : _ans_43_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_43_leadingZeros = _ans_43_leadingZeros_T_93[0] ? 6'h0 : _ans_43_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_43_expRaw_T_1 = 6'h1f - ans_43_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_43_expRaw = ans_43_isZero ? 6'h0 : _ans_43_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_43_shiftAmt_T_2 = ans_43_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_43_shiftAmt = ans_43_expRaw > 6'h3 ? _ans_43_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_43_mantissaRaw_T = ans_43_absClipped >> ans_43_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_43_mantissaRaw = _ans_43_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_43_mantissa = ans_43_expRaw >= 6'h3 ? ans_43_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_43_expAdjusted = ans_43_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_43_exp_T_4 = ans_43_expAdjusted > 7'hf ? 4'hf : ans_43_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_43_exp = ans_43_isZero ? 4'h0 : _ans_43_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_43_fp8 = {ans_43_clippedX[31],ans_43_exp,ans_43_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_44 = {24'h0,linear_bias_44}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_44 = tempSum_44 + biasExtended_44; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_44_sign = sum32_44[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_44_absX_T = ~sum32_44; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_44_absX_T_2 = _ans_44_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_44_absX = ans_44_sign ? _ans_44_absX_T_2 : sum32_44; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_44_shiftedX_T_1 = _GEN_10432 - ans_44_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_44_shiftedX_T_3 = ans_44_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_44_shiftedX = ans_44_sign ? _ans_44_shiftedX_T_1 : _ans_44_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_44_scaledX_T_1 = ans_44_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_44_scaledX = _ans_44_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_44_clippedX_T_2 = ans_44_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_44_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_44_clippedX = ans_44_scaledX > 49'h1c0 ? 49'h1c0 : _ans_44_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_44_absClipped_T_1 = ~ans_44_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_44_absClipped_T_3 = _ans_44_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_44_absClipped = ans_44_clippedX[31] ? _ans_44_absClipped_T_3 : ans_44_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_44_isZero = ans_44_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10918 = {{16'd0}, ans_44_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_4 = _GEN_10918 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_6 = {ans_44_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_8 = _ans_44_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_9 = _ans_44_leadingZeros_T_4 | _ans_44_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10919 = {{8'd0}, _ans_44_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_14 = _GEN_10919 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_16 = {_ans_44_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_18 = _ans_44_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_19 = _ans_44_leadingZeros_T_14 | _ans_44_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10920 = {{4'd0}, _ans_44_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_24 = _GEN_10920 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_26 = {_ans_44_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_28 = _ans_44_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_29 = _ans_44_leadingZeros_T_24 | _ans_44_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10921 = {{2'd0}, _ans_44_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_34 = _GEN_10921 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_36 = {_ans_44_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_38 = _ans_44_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_39 = _ans_44_leadingZeros_T_34 | _ans_44_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10922 = {{1'd0}, _ans_44_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_44 = _GEN_10922 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_46 = {_ans_44_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_48 = _ans_44_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_44_leadingZeros_T_49 = _ans_44_leadingZeros_T_44 | _ans_44_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10923 = {{8'd0}, ans_44_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_55 = _GEN_10923 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_57 = {ans_44_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_59 = _ans_44_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_60 = _ans_44_leadingZeros_T_55 | _ans_44_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10924 = {{4'd0}, _ans_44_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_65 = _GEN_10924 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_67 = {_ans_44_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_69 = _ans_44_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_70 = _ans_44_leadingZeros_T_65 | _ans_44_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10925 = {{2'd0}, _ans_44_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_75 = _GEN_10925 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_77 = {_ans_44_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_79 = _ans_44_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_80 = _ans_44_leadingZeros_T_75 | _ans_44_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10926 = {{1'd0}, _ans_44_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_85 = _GEN_10926 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_87 = {_ans_44_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_89 = _ans_44_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_44_leadingZeros_T_90 = _ans_44_leadingZeros_T_85 | _ans_44_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_44_leadingZeros_T_93 = {_ans_44_leadingZeros_T_49,_ans_44_leadingZeros_T_90,ans_44_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_44_leadingZeros_T_143 = _ans_44_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_144 = _ans_44_leadingZeros_T_93[46] ? 6'h2e : _ans_44_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_145 = _ans_44_leadingZeros_T_93[45] ? 6'h2d : _ans_44_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_146 = _ans_44_leadingZeros_T_93[44] ? 6'h2c : _ans_44_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_147 = _ans_44_leadingZeros_T_93[43] ? 6'h2b : _ans_44_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_148 = _ans_44_leadingZeros_T_93[42] ? 6'h2a : _ans_44_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_149 = _ans_44_leadingZeros_T_93[41] ? 6'h29 : _ans_44_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_150 = _ans_44_leadingZeros_T_93[40] ? 6'h28 : _ans_44_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_151 = _ans_44_leadingZeros_T_93[39] ? 6'h27 : _ans_44_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_152 = _ans_44_leadingZeros_T_93[38] ? 6'h26 : _ans_44_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_153 = _ans_44_leadingZeros_T_93[37] ? 6'h25 : _ans_44_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_154 = _ans_44_leadingZeros_T_93[36] ? 6'h24 : _ans_44_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_155 = _ans_44_leadingZeros_T_93[35] ? 6'h23 : _ans_44_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_156 = _ans_44_leadingZeros_T_93[34] ? 6'h22 : _ans_44_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_157 = _ans_44_leadingZeros_T_93[33] ? 6'h21 : _ans_44_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_158 = _ans_44_leadingZeros_T_93[32] ? 6'h20 : _ans_44_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_159 = _ans_44_leadingZeros_T_93[31] ? 6'h1f : _ans_44_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_160 = _ans_44_leadingZeros_T_93[30] ? 6'h1e : _ans_44_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_161 = _ans_44_leadingZeros_T_93[29] ? 6'h1d : _ans_44_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_162 = _ans_44_leadingZeros_T_93[28] ? 6'h1c : _ans_44_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_163 = _ans_44_leadingZeros_T_93[27] ? 6'h1b : _ans_44_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_164 = _ans_44_leadingZeros_T_93[26] ? 6'h1a : _ans_44_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_165 = _ans_44_leadingZeros_T_93[25] ? 6'h19 : _ans_44_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_166 = _ans_44_leadingZeros_T_93[24] ? 6'h18 : _ans_44_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_167 = _ans_44_leadingZeros_T_93[23] ? 6'h17 : _ans_44_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_168 = _ans_44_leadingZeros_T_93[22] ? 6'h16 : _ans_44_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_169 = _ans_44_leadingZeros_T_93[21] ? 6'h15 : _ans_44_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_170 = _ans_44_leadingZeros_T_93[20] ? 6'h14 : _ans_44_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_171 = _ans_44_leadingZeros_T_93[19] ? 6'h13 : _ans_44_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_172 = _ans_44_leadingZeros_T_93[18] ? 6'h12 : _ans_44_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_173 = _ans_44_leadingZeros_T_93[17] ? 6'h11 : _ans_44_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_174 = _ans_44_leadingZeros_T_93[16] ? 6'h10 : _ans_44_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_175 = _ans_44_leadingZeros_T_93[15] ? 6'hf : _ans_44_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_176 = _ans_44_leadingZeros_T_93[14] ? 6'he : _ans_44_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_177 = _ans_44_leadingZeros_T_93[13] ? 6'hd : _ans_44_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_178 = _ans_44_leadingZeros_T_93[12] ? 6'hc : _ans_44_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_179 = _ans_44_leadingZeros_T_93[11] ? 6'hb : _ans_44_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_180 = _ans_44_leadingZeros_T_93[10] ? 6'ha : _ans_44_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_181 = _ans_44_leadingZeros_T_93[9] ? 6'h9 : _ans_44_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_182 = _ans_44_leadingZeros_T_93[8] ? 6'h8 : _ans_44_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_183 = _ans_44_leadingZeros_T_93[7] ? 6'h7 : _ans_44_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_184 = _ans_44_leadingZeros_T_93[6] ? 6'h6 : _ans_44_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_185 = _ans_44_leadingZeros_T_93[5] ? 6'h5 : _ans_44_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_186 = _ans_44_leadingZeros_T_93[4] ? 6'h4 : _ans_44_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_187 = _ans_44_leadingZeros_T_93[3] ? 6'h3 : _ans_44_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_188 = _ans_44_leadingZeros_T_93[2] ? 6'h2 : _ans_44_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_leadingZeros_T_189 = _ans_44_leadingZeros_T_93[1] ? 6'h1 : _ans_44_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_44_leadingZeros = _ans_44_leadingZeros_T_93[0] ? 6'h0 : _ans_44_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_44_expRaw_T_1 = 6'h1f - ans_44_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_44_expRaw = ans_44_isZero ? 6'h0 : _ans_44_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_44_shiftAmt_T_2 = ans_44_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_44_shiftAmt = ans_44_expRaw > 6'h3 ? _ans_44_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_44_mantissaRaw_T = ans_44_absClipped >> ans_44_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_44_mantissaRaw = _ans_44_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_44_mantissa = ans_44_expRaw >= 6'h3 ? ans_44_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_44_expAdjusted = ans_44_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_44_exp_T_4 = ans_44_expAdjusted > 7'hf ? 4'hf : ans_44_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_44_exp = ans_44_isZero ? 4'h0 : _ans_44_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_44_fp8 = {ans_44_clippedX[31],ans_44_exp,ans_44_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_45 = {24'h0,linear_bias_45}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_45 = tempSum_45 + biasExtended_45; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_45_sign = sum32_45[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_45_absX_T = ~sum32_45; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_45_absX_T_2 = _ans_45_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_45_absX = ans_45_sign ? _ans_45_absX_T_2 : sum32_45; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_45_shiftedX_T_1 = _GEN_10432 - ans_45_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_45_shiftedX_T_3 = ans_45_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_45_shiftedX = ans_45_sign ? _ans_45_shiftedX_T_1 : _ans_45_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_45_scaledX_T_1 = ans_45_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_45_scaledX = _ans_45_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_45_clippedX_T_2 = ans_45_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_45_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_45_clippedX = ans_45_scaledX > 49'h1c0 ? 49'h1c0 : _ans_45_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_45_absClipped_T_1 = ~ans_45_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_45_absClipped_T_3 = _ans_45_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_45_absClipped = ans_45_clippedX[31] ? _ans_45_absClipped_T_3 : ans_45_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_45_isZero = ans_45_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10929 = {{16'd0}, ans_45_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_4 = _GEN_10929 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_6 = {ans_45_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_8 = _ans_45_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_9 = _ans_45_leadingZeros_T_4 | _ans_45_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10930 = {{8'd0}, _ans_45_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_14 = _GEN_10930 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_16 = {_ans_45_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_18 = _ans_45_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_19 = _ans_45_leadingZeros_T_14 | _ans_45_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10931 = {{4'd0}, _ans_45_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_24 = _GEN_10931 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_26 = {_ans_45_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_28 = _ans_45_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_29 = _ans_45_leadingZeros_T_24 | _ans_45_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10932 = {{2'd0}, _ans_45_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_34 = _GEN_10932 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_36 = {_ans_45_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_38 = _ans_45_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_39 = _ans_45_leadingZeros_T_34 | _ans_45_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10933 = {{1'd0}, _ans_45_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_44 = _GEN_10933 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_46 = {_ans_45_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_48 = _ans_45_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_45_leadingZeros_T_49 = _ans_45_leadingZeros_T_44 | _ans_45_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10934 = {{8'd0}, ans_45_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_55 = _GEN_10934 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_57 = {ans_45_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_59 = _ans_45_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_60 = _ans_45_leadingZeros_T_55 | _ans_45_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10935 = {{4'd0}, _ans_45_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_65 = _GEN_10935 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_67 = {_ans_45_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_69 = _ans_45_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_70 = _ans_45_leadingZeros_T_65 | _ans_45_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10936 = {{2'd0}, _ans_45_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_75 = _GEN_10936 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_77 = {_ans_45_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_79 = _ans_45_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_80 = _ans_45_leadingZeros_T_75 | _ans_45_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10937 = {{1'd0}, _ans_45_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_85 = _GEN_10937 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_87 = {_ans_45_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_89 = _ans_45_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_45_leadingZeros_T_90 = _ans_45_leadingZeros_T_85 | _ans_45_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_45_leadingZeros_T_93 = {_ans_45_leadingZeros_T_49,_ans_45_leadingZeros_T_90,ans_45_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_45_leadingZeros_T_143 = _ans_45_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_144 = _ans_45_leadingZeros_T_93[46] ? 6'h2e : _ans_45_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_145 = _ans_45_leadingZeros_T_93[45] ? 6'h2d : _ans_45_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_146 = _ans_45_leadingZeros_T_93[44] ? 6'h2c : _ans_45_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_147 = _ans_45_leadingZeros_T_93[43] ? 6'h2b : _ans_45_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_148 = _ans_45_leadingZeros_T_93[42] ? 6'h2a : _ans_45_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_149 = _ans_45_leadingZeros_T_93[41] ? 6'h29 : _ans_45_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_150 = _ans_45_leadingZeros_T_93[40] ? 6'h28 : _ans_45_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_151 = _ans_45_leadingZeros_T_93[39] ? 6'h27 : _ans_45_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_152 = _ans_45_leadingZeros_T_93[38] ? 6'h26 : _ans_45_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_153 = _ans_45_leadingZeros_T_93[37] ? 6'h25 : _ans_45_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_154 = _ans_45_leadingZeros_T_93[36] ? 6'h24 : _ans_45_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_155 = _ans_45_leadingZeros_T_93[35] ? 6'h23 : _ans_45_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_156 = _ans_45_leadingZeros_T_93[34] ? 6'h22 : _ans_45_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_157 = _ans_45_leadingZeros_T_93[33] ? 6'h21 : _ans_45_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_158 = _ans_45_leadingZeros_T_93[32] ? 6'h20 : _ans_45_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_159 = _ans_45_leadingZeros_T_93[31] ? 6'h1f : _ans_45_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_160 = _ans_45_leadingZeros_T_93[30] ? 6'h1e : _ans_45_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_161 = _ans_45_leadingZeros_T_93[29] ? 6'h1d : _ans_45_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_162 = _ans_45_leadingZeros_T_93[28] ? 6'h1c : _ans_45_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_163 = _ans_45_leadingZeros_T_93[27] ? 6'h1b : _ans_45_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_164 = _ans_45_leadingZeros_T_93[26] ? 6'h1a : _ans_45_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_165 = _ans_45_leadingZeros_T_93[25] ? 6'h19 : _ans_45_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_166 = _ans_45_leadingZeros_T_93[24] ? 6'h18 : _ans_45_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_167 = _ans_45_leadingZeros_T_93[23] ? 6'h17 : _ans_45_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_168 = _ans_45_leadingZeros_T_93[22] ? 6'h16 : _ans_45_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_169 = _ans_45_leadingZeros_T_93[21] ? 6'h15 : _ans_45_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_170 = _ans_45_leadingZeros_T_93[20] ? 6'h14 : _ans_45_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_171 = _ans_45_leadingZeros_T_93[19] ? 6'h13 : _ans_45_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_172 = _ans_45_leadingZeros_T_93[18] ? 6'h12 : _ans_45_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_173 = _ans_45_leadingZeros_T_93[17] ? 6'h11 : _ans_45_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_174 = _ans_45_leadingZeros_T_93[16] ? 6'h10 : _ans_45_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_175 = _ans_45_leadingZeros_T_93[15] ? 6'hf : _ans_45_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_176 = _ans_45_leadingZeros_T_93[14] ? 6'he : _ans_45_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_177 = _ans_45_leadingZeros_T_93[13] ? 6'hd : _ans_45_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_178 = _ans_45_leadingZeros_T_93[12] ? 6'hc : _ans_45_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_179 = _ans_45_leadingZeros_T_93[11] ? 6'hb : _ans_45_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_180 = _ans_45_leadingZeros_T_93[10] ? 6'ha : _ans_45_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_181 = _ans_45_leadingZeros_T_93[9] ? 6'h9 : _ans_45_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_182 = _ans_45_leadingZeros_T_93[8] ? 6'h8 : _ans_45_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_183 = _ans_45_leadingZeros_T_93[7] ? 6'h7 : _ans_45_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_184 = _ans_45_leadingZeros_T_93[6] ? 6'h6 : _ans_45_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_185 = _ans_45_leadingZeros_T_93[5] ? 6'h5 : _ans_45_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_186 = _ans_45_leadingZeros_T_93[4] ? 6'h4 : _ans_45_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_187 = _ans_45_leadingZeros_T_93[3] ? 6'h3 : _ans_45_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_188 = _ans_45_leadingZeros_T_93[2] ? 6'h2 : _ans_45_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_leadingZeros_T_189 = _ans_45_leadingZeros_T_93[1] ? 6'h1 : _ans_45_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_45_leadingZeros = _ans_45_leadingZeros_T_93[0] ? 6'h0 : _ans_45_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_45_expRaw_T_1 = 6'h1f - ans_45_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_45_expRaw = ans_45_isZero ? 6'h0 : _ans_45_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_45_shiftAmt_T_2 = ans_45_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_45_shiftAmt = ans_45_expRaw > 6'h3 ? _ans_45_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_45_mantissaRaw_T = ans_45_absClipped >> ans_45_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_45_mantissaRaw = _ans_45_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_45_mantissa = ans_45_expRaw >= 6'h3 ? ans_45_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_45_expAdjusted = ans_45_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_45_exp_T_4 = ans_45_expAdjusted > 7'hf ? 4'hf : ans_45_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_45_exp = ans_45_isZero ? 4'h0 : _ans_45_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_45_fp8 = {ans_45_clippedX[31],ans_45_exp,ans_45_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_46 = {24'h0,linear_bias_46}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_46 = tempSum_46 + biasExtended_46; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_46_sign = sum32_46[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_46_absX_T = ~sum32_46; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_46_absX_T_2 = _ans_46_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_46_absX = ans_46_sign ? _ans_46_absX_T_2 : sum32_46; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_46_shiftedX_T_1 = _GEN_10432 - ans_46_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_46_shiftedX_T_3 = ans_46_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_46_shiftedX = ans_46_sign ? _ans_46_shiftedX_T_1 : _ans_46_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_46_scaledX_T_1 = ans_46_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_46_scaledX = _ans_46_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_46_clippedX_T_2 = ans_46_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_46_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_46_clippedX = ans_46_scaledX > 49'h1c0 ? 49'h1c0 : _ans_46_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_46_absClipped_T_1 = ~ans_46_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_46_absClipped_T_3 = _ans_46_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_46_absClipped = ans_46_clippedX[31] ? _ans_46_absClipped_T_3 : ans_46_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_46_isZero = ans_46_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10940 = {{16'd0}, ans_46_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_4 = _GEN_10940 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_6 = {ans_46_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_8 = _ans_46_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_9 = _ans_46_leadingZeros_T_4 | _ans_46_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10941 = {{8'd0}, _ans_46_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_14 = _GEN_10941 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_16 = {_ans_46_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_18 = _ans_46_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_19 = _ans_46_leadingZeros_T_14 | _ans_46_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10942 = {{4'd0}, _ans_46_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_24 = _GEN_10942 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_26 = {_ans_46_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_28 = _ans_46_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_29 = _ans_46_leadingZeros_T_24 | _ans_46_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10943 = {{2'd0}, _ans_46_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_34 = _GEN_10943 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_36 = {_ans_46_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_38 = _ans_46_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_39 = _ans_46_leadingZeros_T_34 | _ans_46_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10944 = {{1'd0}, _ans_46_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_44 = _GEN_10944 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_46 = {_ans_46_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_48 = _ans_46_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_46_leadingZeros_T_49 = _ans_46_leadingZeros_T_44 | _ans_46_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10945 = {{8'd0}, ans_46_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_55 = _GEN_10945 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_57 = {ans_46_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_59 = _ans_46_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_60 = _ans_46_leadingZeros_T_55 | _ans_46_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10946 = {{4'd0}, _ans_46_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_65 = _GEN_10946 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_67 = {_ans_46_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_69 = _ans_46_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_70 = _ans_46_leadingZeros_T_65 | _ans_46_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10947 = {{2'd0}, _ans_46_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_75 = _GEN_10947 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_77 = {_ans_46_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_79 = _ans_46_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_80 = _ans_46_leadingZeros_T_75 | _ans_46_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10948 = {{1'd0}, _ans_46_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_85 = _GEN_10948 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_87 = {_ans_46_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_89 = _ans_46_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_46_leadingZeros_T_90 = _ans_46_leadingZeros_T_85 | _ans_46_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_46_leadingZeros_T_93 = {_ans_46_leadingZeros_T_49,_ans_46_leadingZeros_T_90,ans_46_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_46_leadingZeros_T_143 = _ans_46_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_144 = _ans_46_leadingZeros_T_93[46] ? 6'h2e : _ans_46_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_145 = _ans_46_leadingZeros_T_93[45] ? 6'h2d : _ans_46_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_146 = _ans_46_leadingZeros_T_93[44] ? 6'h2c : _ans_46_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_147 = _ans_46_leadingZeros_T_93[43] ? 6'h2b : _ans_46_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_148 = _ans_46_leadingZeros_T_93[42] ? 6'h2a : _ans_46_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_149 = _ans_46_leadingZeros_T_93[41] ? 6'h29 : _ans_46_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_150 = _ans_46_leadingZeros_T_93[40] ? 6'h28 : _ans_46_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_151 = _ans_46_leadingZeros_T_93[39] ? 6'h27 : _ans_46_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_152 = _ans_46_leadingZeros_T_93[38] ? 6'h26 : _ans_46_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_153 = _ans_46_leadingZeros_T_93[37] ? 6'h25 : _ans_46_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_154 = _ans_46_leadingZeros_T_93[36] ? 6'h24 : _ans_46_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_155 = _ans_46_leadingZeros_T_93[35] ? 6'h23 : _ans_46_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_156 = _ans_46_leadingZeros_T_93[34] ? 6'h22 : _ans_46_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_157 = _ans_46_leadingZeros_T_93[33] ? 6'h21 : _ans_46_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_158 = _ans_46_leadingZeros_T_93[32] ? 6'h20 : _ans_46_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_159 = _ans_46_leadingZeros_T_93[31] ? 6'h1f : _ans_46_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_160 = _ans_46_leadingZeros_T_93[30] ? 6'h1e : _ans_46_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_161 = _ans_46_leadingZeros_T_93[29] ? 6'h1d : _ans_46_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_162 = _ans_46_leadingZeros_T_93[28] ? 6'h1c : _ans_46_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_163 = _ans_46_leadingZeros_T_93[27] ? 6'h1b : _ans_46_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_164 = _ans_46_leadingZeros_T_93[26] ? 6'h1a : _ans_46_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_165 = _ans_46_leadingZeros_T_93[25] ? 6'h19 : _ans_46_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_166 = _ans_46_leadingZeros_T_93[24] ? 6'h18 : _ans_46_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_167 = _ans_46_leadingZeros_T_93[23] ? 6'h17 : _ans_46_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_168 = _ans_46_leadingZeros_T_93[22] ? 6'h16 : _ans_46_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_169 = _ans_46_leadingZeros_T_93[21] ? 6'h15 : _ans_46_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_170 = _ans_46_leadingZeros_T_93[20] ? 6'h14 : _ans_46_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_171 = _ans_46_leadingZeros_T_93[19] ? 6'h13 : _ans_46_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_172 = _ans_46_leadingZeros_T_93[18] ? 6'h12 : _ans_46_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_173 = _ans_46_leadingZeros_T_93[17] ? 6'h11 : _ans_46_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_174 = _ans_46_leadingZeros_T_93[16] ? 6'h10 : _ans_46_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_175 = _ans_46_leadingZeros_T_93[15] ? 6'hf : _ans_46_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_176 = _ans_46_leadingZeros_T_93[14] ? 6'he : _ans_46_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_177 = _ans_46_leadingZeros_T_93[13] ? 6'hd : _ans_46_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_178 = _ans_46_leadingZeros_T_93[12] ? 6'hc : _ans_46_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_179 = _ans_46_leadingZeros_T_93[11] ? 6'hb : _ans_46_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_180 = _ans_46_leadingZeros_T_93[10] ? 6'ha : _ans_46_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_181 = _ans_46_leadingZeros_T_93[9] ? 6'h9 : _ans_46_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_182 = _ans_46_leadingZeros_T_93[8] ? 6'h8 : _ans_46_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_183 = _ans_46_leadingZeros_T_93[7] ? 6'h7 : _ans_46_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_184 = _ans_46_leadingZeros_T_93[6] ? 6'h6 : _ans_46_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_185 = _ans_46_leadingZeros_T_93[5] ? 6'h5 : _ans_46_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_186 = _ans_46_leadingZeros_T_93[4] ? 6'h4 : _ans_46_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_187 = _ans_46_leadingZeros_T_93[3] ? 6'h3 : _ans_46_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_188 = _ans_46_leadingZeros_T_93[2] ? 6'h2 : _ans_46_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_leadingZeros_T_189 = _ans_46_leadingZeros_T_93[1] ? 6'h1 : _ans_46_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_46_leadingZeros = _ans_46_leadingZeros_T_93[0] ? 6'h0 : _ans_46_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_46_expRaw_T_1 = 6'h1f - ans_46_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_46_expRaw = ans_46_isZero ? 6'h0 : _ans_46_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_46_shiftAmt_T_2 = ans_46_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_46_shiftAmt = ans_46_expRaw > 6'h3 ? _ans_46_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_46_mantissaRaw_T = ans_46_absClipped >> ans_46_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_46_mantissaRaw = _ans_46_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_46_mantissa = ans_46_expRaw >= 6'h3 ? ans_46_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_46_expAdjusted = ans_46_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_46_exp_T_4 = ans_46_expAdjusted > 7'hf ? 4'hf : ans_46_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_46_exp = ans_46_isZero ? 4'h0 : _ans_46_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_46_fp8 = {ans_46_clippedX[31],ans_46_exp,ans_46_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_47 = {24'h0,linear_bias_47}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_47 = tempSum_47 + biasExtended_47; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_47_sign = sum32_47[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_47_absX_T = ~sum32_47; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_47_absX_T_2 = _ans_47_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_47_absX = ans_47_sign ? _ans_47_absX_T_2 : sum32_47; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_47_shiftedX_T_1 = _GEN_10432 - ans_47_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_47_shiftedX_T_3 = ans_47_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_47_shiftedX = ans_47_sign ? _ans_47_shiftedX_T_1 : _ans_47_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_47_scaledX_T_1 = ans_47_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_47_scaledX = _ans_47_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_47_clippedX_T_2 = ans_47_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_47_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_47_clippedX = ans_47_scaledX > 49'h1c0 ? 49'h1c0 : _ans_47_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_47_absClipped_T_1 = ~ans_47_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_47_absClipped_T_3 = _ans_47_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_47_absClipped = ans_47_clippedX[31] ? _ans_47_absClipped_T_3 : ans_47_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_47_isZero = ans_47_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10951 = {{16'd0}, ans_47_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_4 = _GEN_10951 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_6 = {ans_47_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_8 = _ans_47_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_9 = _ans_47_leadingZeros_T_4 | _ans_47_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10952 = {{8'd0}, _ans_47_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_14 = _GEN_10952 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_16 = {_ans_47_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_18 = _ans_47_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_19 = _ans_47_leadingZeros_T_14 | _ans_47_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10953 = {{4'd0}, _ans_47_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_24 = _GEN_10953 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_26 = {_ans_47_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_28 = _ans_47_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_29 = _ans_47_leadingZeros_T_24 | _ans_47_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10954 = {{2'd0}, _ans_47_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_34 = _GEN_10954 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_36 = {_ans_47_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_38 = _ans_47_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_39 = _ans_47_leadingZeros_T_34 | _ans_47_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10955 = {{1'd0}, _ans_47_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_44 = _GEN_10955 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_46 = {_ans_47_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_48 = _ans_47_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_47_leadingZeros_T_49 = _ans_47_leadingZeros_T_44 | _ans_47_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10956 = {{8'd0}, ans_47_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_55 = _GEN_10956 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_57 = {ans_47_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_59 = _ans_47_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_60 = _ans_47_leadingZeros_T_55 | _ans_47_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10957 = {{4'd0}, _ans_47_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_65 = _GEN_10957 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_67 = {_ans_47_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_69 = _ans_47_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_70 = _ans_47_leadingZeros_T_65 | _ans_47_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10958 = {{2'd0}, _ans_47_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_75 = _GEN_10958 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_77 = {_ans_47_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_79 = _ans_47_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_80 = _ans_47_leadingZeros_T_75 | _ans_47_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10959 = {{1'd0}, _ans_47_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_85 = _GEN_10959 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_87 = {_ans_47_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_89 = _ans_47_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_47_leadingZeros_T_90 = _ans_47_leadingZeros_T_85 | _ans_47_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_47_leadingZeros_T_93 = {_ans_47_leadingZeros_T_49,_ans_47_leadingZeros_T_90,ans_47_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_47_leadingZeros_T_143 = _ans_47_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_144 = _ans_47_leadingZeros_T_93[46] ? 6'h2e : _ans_47_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_145 = _ans_47_leadingZeros_T_93[45] ? 6'h2d : _ans_47_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_146 = _ans_47_leadingZeros_T_93[44] ? 6'h2c : _ans_47_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_147 = _ans_47_leadingZeros_T_93[43] ? 6'h2b : _ans_47_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_148 = _ans_47_leadingZeros_T_93[42] ? 6'h2a : _ans_47_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_149 = _ans_47_leadingZeros_T_93[41] ? 6'h29 : _ans_47_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_150 = _ans_47_leadingZeros_T_93[40] ? 6'h28 : _ans_47_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_151 = _ans_47_leadingZeros_T_93[39] ? 6'h27 : _ans_47_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_152 = _ans_47_leadingZeros_T_93[38] ? 6'h26 : _ans_47_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_153 = _ans_47_leadingZeros_T_93[37] ? 6'h25 : _ans_47_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_154 = _ans_47_leadingZeros_T_93[36] ? 6'h24 : _ans_47_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_155 = _ans_47_leadingZeros_T_93[35] ? 6'h23 : _ans_47_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_156 = _ans_47_leadingZeros_T_93[34] ? 6'h22 : _ans_47_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_157 = _ans_47_leadingZeros_T_93[33] ? 6'h21 : _ans_47_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_158 = _ans_47_leadingZeros_T_93[32] ? 6'h20 : _ans_47_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_159 = _ans_47_leadingZeros_T_93[31] ? 6'h1f : _ans_47_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_160 = _ans_47_leadingZeros_T_93[30] ? 6'h1e : _ans_47_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_161 = _ans_47_leadingZeros_T_93[29] ? 6'h1d : _ans_47_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_162 = _ans_47_leadingZeros_T_93[28] ? 6'h1c : _ans_47_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_163 = _ans_47_leadingZeros_T_93[27] ? 6'h1b : _ans_47_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_164 = _ans_47_leadingZeros_T_93[26] ? 6'h1a : _ans_47_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_165 = _ans_47_leadingZeros_T_93[25] ? 6'h19 : _ans_47_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_166 = _ans_47_leadingZeros_T_93[24] ? 6'h18 : _ans_47_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_167 = _ans_47_leadingZeros_T_93[23] ? 6'h17 : _ans_47_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_168 = _ans_47_leadingZeros_T_93[22] ? 6'h16 : _ans_47_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_169 = _ans_47_leadingZeros_T_93[21] ? 6'h15 : _ans_47_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_170 = _ans_47_leadingZeros_T_93[20] ? 6'h14 : _ans_47_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_171 = _ans_47_leadingZeros_T_93[19] ? 6'h13 : _ans_47_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_172 = _ans_47_leadingZeros_T_93[18] ? 6'h12 : _ans_47_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_173 = _ans_47_leadingZeros_T_93[17] ? 6'h11 : _ans_47_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_174 = _ans_47_leadingZeros_T_93[16] ? 6'h10 : _ans_47_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_175 = _ans_47_leadingZeros_T_93[15] ? 6'hf : _ans_47_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_176 = _ans_47_leadingZeros_T_93[14] ? 6'he : _ans_47_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_177 = _ans_47_leadingZeros_T_93[13] ? 6'hd : _ans_47_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_178 = _ans_47_leadingZeros_T_93[12] ? 6'hc : _ans_47_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_179 = _ans_47_leadingZeros_T_93[11] ? 6'hb : _ans_47_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_180 = _ans_47_leadingZeros_T_93[10] ? 6'ha : _ans_47_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_181 = _ans_47_leadingZeros_T_93[9] ? 6'h9 : _ans_47_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_182 = _ans_47_leadingZeros_T_93[8] ? 6'h8 : _ans_47_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_183 = _ans_47_leadingZeros_T_93[7] ? 6'h7 : _ans_47_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_184 = _ans_47_leadingZeros_T_93[6] ? 6'h6 : _ans_47_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_185 = _ans_47_leadingZeros_T_93[5] ? 6'h5 : _ans_47_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_186 = _ans_47_leadingZeros_T_93[4] ? 6'h4 : _ans_47_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_187 = _ans_47_leadingZeros_T_93[3] ? 6'h3 : _ans_47_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_188 = _ans_47_leadingZeros_T_93[2] ? 6'h2 : _ans_47_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_leadingZeros_T_189 = _ans_47_leadingZeros_T_93[1] ? 6'h1 : _ans_47_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_47_leadingZeros = _ans_47_leadingZeros_T_93[0] ? 6'h0 : _ans_47_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_47_expRaw_T_1 = 6'h1f - ans_47_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_47_expRaw = ans_47_isZero ? 6'h0 : _ans_47_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_47_shiftAmt_T_2 = ans_47_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_47_shiftAmt = ans_47_expRaw > 6'h3 ? _ans_47_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_47_mantissaRaw_T = ans_47_absClipped >> ans_47_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_47_mantissaRaw = _ans_47_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_47_mantissa = ans_47_expRaw >= 6'h3 ? ans_47_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_47_expAdjusted = ans_47_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_47_exp_T_4 = ans_47_expAdjusted > 7'hf ? 4'hf : ans_47_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_47_exp = ans_47_isZero ? 4'h0 : _ans_47_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_47_fp8 = {ans_47_clippedX[31],ans_47_exp,ans_47_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_48 = {24'h0,linear_bias_48}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_48 = tempSum_48 + biasExtended_48; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_48_sign = sum32_48[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_48_absX_T = ~sum32_48; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_48_absX_T_2 = _ans_48_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_48_absX = ans_48_sign ? _ans_48_absX_T_2 : sum32_48; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_48_shiftedX_T_1 = _GEN_10432 - ans_48_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_48_shiftedX_T_3 = ans_48_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_48_shiftedX = ans_48_sign ? _ans_48_shiftedX_T_1 : _ans_48_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_48_scaledX_T_1 = ans_48_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_48_scaledX = _ans_48_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_48_clippedX_T_2 = ans_48_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_48_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_48_clippedX = ans_48_scaledX > 49'h1c0 ? 49'h1c0 : _ans_48_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_48_absClipped_T_1 = ~ans_48_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_48_absClipped_T_3 = _ans_48_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_48_absClipped = ans_48_clippedX[31] ? _ans_48_absClipped_T_3 : ans_48_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_48_isZero = ans_48_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10962 = {{16'd0}, ans_48_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_4 = _GEN_10962 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_6 = {ans_48_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_8 = _ans_48_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_9 = _ans_48_leadingZeros_T_4 | _ans_48_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10963 = {{8'd0}, _ans_48_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_14 = _GEN_10963 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_16 = {_ans_48_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_18 = _ans_48_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_19 = _ans_48_leadingZeros_T_14 | _ans_48_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10964 = {{4'd0}, _ans_48_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_24 = _GEN_10964 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_26 = {_ans_48_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_28 = _ans_48_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_29 = _ans_48_leadingZeros_T_24 | _ans_48_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10965 = {{2'd0}, _ans_48_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_34 = _GEN_10965 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_36 = {_ans_48_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_38 = _ans_48_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_39 = _ans_48_leadingZeros_T_34 | _ans_48_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10966 = {{1'd0}, _ans_48_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_44 = _GEN_10966 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_46 = {_ans_48_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_48 = _ans_48_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_48_leadingZeros_T_49 = _ans_48_leadingZeros_T_44 | _ans_48_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10967 = {{8'd0}, ans_48_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_55 = _GEN_10967 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_57 = {ans_48_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_59 = _ans_48_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_60 = _ans_48_leadingZeros_T_55 | _ans_48_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10968 = {{4'd0}, _ans_48_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_65 = _GEN_10968 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_67 = {_ans_48_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_69 = _ans_48_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_70 = _ans_48_leadingZeros_T_65 | _ans_48_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10969 = {{2'd0}, _ans_48_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_75 = _GEN_10969 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_77 = {_ans_48_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_79 = _ans_48_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_80 = _ans_48_leadingZeros_T_75 | _ans_48_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10970 = {{1'd0}, _ans_48_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_85 = _GEN_10970 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_87 = {_ans_48_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_89 = _ans_48_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_48_leadingZeros_T_90 = _ans_48_leadingZeros_T_85 | _ans_48_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_48_leadingZeros_T_93 = {_ans_48_leadingZeros_T_49,_ans_48_leadingZeros_T_90,ans_48_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_48_leadingZeros_T_143 = _ans_48_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_144 = _ans_48_leadingZeros_T_93[46] ? 6'h2e : _ans_48_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_145 = _ans_48_leadingZeros_T_93[45] ? 6'h2d : _ans_48_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_146 = _ans_48_leadingZeros_T_93[44] ? 6'h2c : _ans_48_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_147 = _ans_48_leadingZeros_T_93[43] ? 6'h2b : _ans_48_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_148 = _ans_48_leadingZeros_T_93[42] ? 6'h2a : _ans_48_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_149 = _ans_48_leadingZeros_T_93[41] ? 6'h29 : _ans_48_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_150 = _ans_48_leadingZeros_T_93[40] ? 6'h28 : _ans_48_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_151 = _ans_48_leadingZeros_T_93[39] ? 6'h27 : _ans_48_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_152 = _ans_48_leadingZeros_T_93[38] ? 6'h26 : _ans_48_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_153 = _ans_48_leadingZeros_T_93[37] ? 6'h25 : _ans_48_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_154 = _ans_48_leadingZeros_T_93[36] ? 6'h24 : _ans_48_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_155 = _ans_48_leadingZeros_T_93[35] ? 6'h23 : _ans_48_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_156 = _ans_48_leadingZeros_T_93[34] ? 6'h22 : _ans_48_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_157 = _ans_48_leadingZeros_T_93[33] ? 6'h21 : _ans_48_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_158 = _ans_48_leadingZeros_T_93[32] ? 6'h20 : _ans_48_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_159 = _ans_48_leadingZeros_T_93[31] ? 6'h1f : _ans_48_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_160 = _ans_48_leadingZeros_T_93[30] ? 6'h1e : _ans_48_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_161 = _ans_48_leadingZeros_T_93[29] ? 6'h1d : _ans_48_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_162 = _ans_48_leadingZeros_T_93[28] ? 6'h1c : _ans_48_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_163 = _ans_48_leadingZeros_T_93[27] ? 6'h1b : _ans_48_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_164 = _ans_48_leadingZeros_T_93[26] ? 6'h1a : _ans_48_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_165 = _ans_48_leadingZeros_T_93[25] ? 6'h19 : _ans_48_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_166 = _ans_48_leadingZeros_T_93[24] ? 6'h18 : _ans_48_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_167 = _ans_48_leadingZeros_T_93[23] ? 6'h17 : _ans_48_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_168 = _ans_48_leadingZeros_T_93[22] ? 6'h16 : _ans_48_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_169 = _ans_48_leadingZeros_T_93[21] ? 6'h15 : _ans_48_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_170 = _ans_48_leadingZeros_T_93[20] ? 6'h14 : _ans_48_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_171 = _ans_48_leadingZeros_T_93[19] ? 6'h13 : _ans_48_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_172 = _ans_48_leadingZeros_T_93[18] ? 6'h12 : _ans_48_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_173 = _ans_48_leadingZeros_T_93[17] ? 6'h11 : _ans_48_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_174 = _ans_48_leadingZeros_T_93[16] ? 6'h10 : _ans_48_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_175 = _ans_48_leadingZeros_T_93[15] ? 6'hf : _ans_48_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_176 = _ans_48_leadingZeros_T_93[14] ? 6'he : _ans_48_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_177 = _ans_48_leadingZeros_T_93[13] ? 6'hd : _ans_48_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_178 = _ans_48_leadingZeros_T_93[12] ? 6'hc : _ans_48_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_179 = _ans_48_leadingZeros_T_93[11] ? 6'hb : _ans_48_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_180 = _ans_48_leadingZeros_T_93[10] ? 6'ha : _ans_48_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_181 = _ans_48_leadingZeros_T_93[9] ? 6'h9 : _ans_48_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_182 = _ans_48_leadingZeros_T_93[8] ? 6'h8 : _ans_48_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_183 = _ans_48_leadingZeros_T_93[7] ? 6'h7 : _ans_48_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_184 = _ans_48_leadingZeros_T_93[6] ? 6'h6 : _ans_48_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_185 = _ans_48_leadingZeros_T_93[5] ? 6'h5 : _ans_48_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_186 = _ans_48_leadingZeros_T_93[4] ? 6'h4 : _ans_48_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_187 = _ans_48_leadingZeros_T_93[3] ? 6'h3 : _ans_48_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_188 = _ans_48_leadingZeros_T_93[2] ? 6'h2 : _ans_48_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_leadingZeros_T_189 = _ans_48_leadingZeros_T_93[1] ? 6'h1 : _ans_48_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_48_leadingZeros = _ans_48_leadingZeros_T_93[0] ? 6'h0 : _ans_48_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_48_expRaw_T_1 = 6'h1f - ans_48_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_48_expRaw = ans_48_isZero ? 6'h0 : _ans_48_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_48_shiftAmt_T_2 = ans_48_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_48_shiftAmt = ans_48_expRaw > 6'h3 ? _ans_48_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_48_mantissaRaw_T = ans_48_absClipped >> ans_48_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_48_mantissaRaw = _ans_48_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_48_mantissa = ans_48_expRaw >= 6'h3 ? ans_48_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_48_expAdjusted = ans_48_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_48_exp_T_4 = ans_48_expAdjusted > 7'hf ? 4'hf : ans_48_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_48_exp = ans_48_isZero ? 4'h0 : _ans_48_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_48_fp8 = {ans_48_clippedX[31],ans_48_exp,ans_48_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_49 = {24'h0,linear_bias_49}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_49 = tempSum_49 + biasExtended_49; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_49_sign = sum32_49[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_49_absX_T = ~sum32_49; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_49_absX_T_2 = _ans_49_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_49_absX = ans_49_sign ? _ans_49_absX_T_2 : sum32_49; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_49_shiftedX_T_1 = _GEN_10432 - ans_49_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_49_shiftedX_T_3 = ans_49_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_49_shiftedX = ans_49_sign ? _ans_49_shiftedX_T_1 : _ans_49_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_49_scaledX_T_1 = ans_49_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_49_scaledX = _ans_49_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_49_clippedX_T_2 = ans_49_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_49_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_49_clippedX = ans_49_scaledX > 49'h1c0 ? 49'h1c0 : _ans_49_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_49_absClipped_T_1 = ~ans_49_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_49_absClipped_T_3 = _ans_49_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_49_absClipped = ans_49_clippedX[31] ? _ans_49_absClipped_T_3 : ans_49_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_49_isZero = ans_49_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10973 = {{16'd0}, ans_49_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_4 = _GEN_10973 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_6 = {ans_49_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_8 = _ans_49_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_9 = _ans_49_leadingZeros_T_4 | _ans_49_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10974 = {{8'd0}, _ans_49_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_14 = _GEN_10974 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_16 = {_ans_49_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_18 = _ans_49_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_19 = _ans_49_leadingZeros_T_14 | _ans_49_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10975 = {{4'd0}, _ans_49_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_24 = _GEN_10975 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_26 = {_ans_49_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_28 = _ans_49_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_29 = _ans_49_leadingZeros_T_24 | _ans_49_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10976 = {{2'd0}, _ans_49_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_34 = _GEN_10976 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_36 = {_ans_49_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_38 = _ans_49_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_39 = _ans_49_leadingZeros_T_34 | _ans_49_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10977 = {{1'd0}, _ans_49_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_44 = _GEN_10977 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_46 = {_ans_49_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_48 = _ans_49_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_49_leadingZeros_T_49 = _ans_49_leadingZeros_T_44 | _ans_49_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10978 = {{8'd0}, ans_49_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_55 = _GEN_10978 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_57 = {ans_49_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_59 = _ans_49_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_60 = _ans_49_leadingZeros_T_55 | _ans_49_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10979 = {{4'd0}, _ans_49_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_65 = _GEN_10979 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_67 = {_ans_49_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_69 = _ans_49_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_70 = _ans_49_leadingZeros_T_65 | _ans_49_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10980 = {{2'd0}, _ans_49_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_75 = _GEN_10980 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_77 = {_ans_49_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_79 = _ans_49_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_80 = _ans_49_leadingZeros_T_75 | _ans_49_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10981 = {{1'd0}, _ans_49_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_85 = _GEN_10981 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_87 = {_ans_49_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_89 = _ans_49_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_49_leadingZeros_T_90 = _ans_49_leadingZeros_T_85 | _ans_49_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_49_leadingZeros_T_93 = {_ans_49_leadingZeros_T_49,_ans_49_leadingZeros_T_90,ans_49_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_49_leadingZeros_T_143 = _ans_49_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_144 = _ans_49_leadingZeros_T_93[46] ? 6'h2e : _ans_49_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_145 = _ans_49_leadingZeros_T_93[45] ? 6'h2d : _ans_49_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_146 = _ans_49_leadingZeros_T_93[44] ? 6'h2c : _ans_49_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_147 = _ans_49_leadingZeros_T_93[43] ? 6'h2b : _ans_49_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_148 = _ans_49_leadingZeros_T_93[42] ? 6'h2a : _ans_49_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_149 = _ans_49_leadingZeros_T_93[41] ? 6'h29 : _ans_49_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_150 = _ans_49_leadingZeros_T_93[40] ? 6'h28 : _ans_49_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_151 = _ans_49_leadingZeros_T_93[39] ? 6'h27 : _ans_49_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_152 = _ans_49_leadingZeros_T_93[38] ? 6'h26 : _ans_49_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_153 = _ans_49_leadingZeros_T_93[37] ? 6'h25 : _ans_49_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_154 = _ans_49_leadingZeros_T_93[36] ? 6'h24 : _ans_49_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_155 = _ans_49_leadingZeros_T_93[35] ? 6'h23 : _ans_49_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_156 = _ans_49_leadingZeros_T_93[34] ? 6'h22 : _ans_49_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_157 = _ans_49_leadingZeros_T_93[33] ? 6'h21 : _ans_49_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_158 = _ans_49_leadingZeros_T_93[32] ? 6'h20 : _ans_49_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_159 = _ans_49_leadingZeros_T_93[31] ? 6'h1f : _ans_49_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_160 = _ans_49_leadingZeros_T_93[30] ? 6'h1e : _ans_49_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_161 = _ans_49_leadingZeros_T_93[29] ? 6'h1d : _ans_49_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_162 = _ans_49_leadingZeros_T_93[28] ? 6'h1c : _ans_49_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_163 = _ans_49_leadingZeros_T_93[27] ? 6'h1b : _ans_49_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_164 = _ans_49_leadingZeros_T_93[26] ? 6'h1a : _ans_49_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_165 = _ans_49_leadingZeros_T_93[25] ? 6'h19 : _ans_49_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_166 = _ans_49_leadingZeros_T_93[24] ? 6'h18 : _ans_49_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_167 = _ans_49_leadingZeros_T_93[23] ? 6'h17 : _ans_49_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_168 = _ans_49_leadingZeros_T_93[22] ? 6'h16 : _ans_49_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_169 = _ans_49_leadingZeros_T_93[21] ? 6'h15 : _ans_49_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_170 = _ans_49_leadingZeros_T_93[20] ? 6'h14 : _ans_49_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_171 = _ans_49_leadingZeros_T_93[19] ? 6'h13 : _ans_49_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_172 = _ans_49_leadingZeros_T_93[18] ? 6'h12 : _ans_49_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_173 = _ans_49_leadingZeros_T_93[17] ? 6'h11 : _ans_49_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_174 = _ans_49_leadingZeros_T_93[16] ? 6'h10 : _ans_49_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_175 = _ans_49_leadingZeros_T_93[15] ? 6'hf : _ans_49_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_176 = _ans_49_leadingZeros_T_93[14] ? 6'he : _ans_49_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_177 = _ans_49_leadingZeros_T_93[13] ? 6'hd : _ans_49_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_178 = _ans_49_leadingZeros_T_93[12] ? 6'hc : _ans_49_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_179 = _ans_49_leadingZeros_T_93[11] ? 6'hb : _ans_49_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_180 = _ans_49_leadingZeros_T_93[10] ? 6'ha : _ans_49_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_181 = _ans_49_leadingZeros_T_93[9] ? 6'h9 : _ans_49_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_182 = _ans_49_leadingZeros_T_93[8] ? 6'h8 : _ans_49_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_183 = _ans_49_leadingZeros_T_93[7] ? 6'h7 : _ans_49_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_184 = _ans_49_leadingZeros_T_93[6] ? 6'h6 : _ans_49_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_185 = _ans_49_leadingZeros_T_93[5] ? 6'h5 : _ans_49_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_186 = _ans_49_leadingZeros_T_93[4] ? 6'h4 : _ans_49_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_187 = _ans_49_leadingZeros_T_93[3] ? 6'h3 : _ans_49_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_188 = _ans_49_leadingZeros_T_93[2] ? 6'h2 : _ans_49_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_leadingZeros_T_189 = _ans_49_leadingZeros_T_93[1] ? 6'h1 : _ans_49_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_49_leadingZeros = _ans_49_leadingZeros_T_93[0] ? 6'h0 : _ans_49_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_49_expRaw_T_1 = 6'h1f - ans_49_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_49_expRaw = ans_49_isZero ? 6'h0 : _ans_49_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_49_shiftAmt_T_2 = ans_49_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_49_shiftAmt = ans_49_expRaw > 6'h3 ? _ans_49_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_49_mantissaRaw_T = ans_49_absClipped >> ans_49_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_49_mantissaRaw = _ans_49_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_49_mantissa = ans_49_expRaw >= 6'h3 ? ans_49_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_49_expAdjusted = ans_49_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_49_exp_T_4 = ans_49_expAdjusted > 7'hf ? 4'hf : ans_49_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_49_exp = ans_49_isZero ? 4'h0 : _ans_49_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_49_fp8 = {ans_49_clippedX[31],ans_49_exp,ans_49_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_50 = {24'h0,linear_bias_50}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_50 = tempSum_50 + biasExtended_50; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_50_sign = sum32_50[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_50_absX_T = ~sum32_50; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_50_absX_T_2 = _ans_50_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_50_absX = ans_50_sign ? _ans_50_absX_T_2 : sum32_50; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_50_shiftedX_T_1 = _GEN_10432 - ans_50_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_50_shiftedX_T_3 = ans_50_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_50_shiftedX = ans_50_sign ? _ans_50_shiftedX_T_1 : _ans_50_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_50_scaledX_T_1 = ans_50_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_50_scaledX = _ans_50_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_50_clippedX_T_2 = ans_50_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_50_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_50_clippedX = ans_50_scaledX > 49'h1c0 ? 49'h1c0 : _ans_50_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_50_absClipped_T_1 = ~ans_50_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_50_absClipped_T_3 = _ans_50_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_50_absClipped = ans_50_clippedX[31] ? _ans_50_absClipped_T_3 : ans_50_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_50_isZero = ans_50_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10984 = {{16'd0}, ans_50_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_4 = _GEN_10984 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_6 = {ans_50_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_8 = _ans_50_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_9 = _ans_50_leadingZeros_T_4 | _ans_50_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10985 = {{8'd0}, _ans_50_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_14 = _GEN_10985 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_16 = {_ans_50_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_18 = _ans_50_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_19 = _ans_50_leadingZeros_T_14 | _ans_50_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10986 = {{4'd0}, _ans_50_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_24 = _GEN_10986 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_26 = {_ans_50_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_28 = _ans_50_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_29 = _ans_50_leadingZeros_T_24 | _ans_50_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10987 = {{2'd0}, _ans_50_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_34 = _GEN_10987 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_36 = {_ans_50_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_38 = _ans_50_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_39 = _ans_50_leadingZeros_T_34 | _ans_50_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10988 = {{1'd0}, _ans_50_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_44 = _GEN_10988 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_46 = {_ans_50_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_48 = _ans_50_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_50_leadingZeros_T_49 = _ans_50_leadingZeros_T_44 | _ans_50_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10989 = {{8'd0}, ans_50_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_55 = _GEN_10989 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_57 = {ans_50_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_59 = _ans_50_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_60 = _ans_50_leadingZeros_T_55 | _ans_50_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10990 = {{4'd0}, _ans_50_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_65 = _GEN_10990 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_67 = {_ans_50_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_69 = _ans_50_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_70 = _ans_50_leadingZeros_T_65 | _ans_50_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10991 = {{2'd0}, _ans_50_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_75 = _GEN_10991 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_77 = {_ans_50_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_79 = _ans_50_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_80 = _ans_50_leadingZeros_T_75 | _ans_50_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_10992 = {{1'd0}, _ans_50_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_85 = _GEN_10992 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_87 = {_ans_50_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_89 = _ans_50_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_50_leadingZeros_T_90 = _ans_50_leadingZeros_T_85 | _ans_50_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_50_leadingZeros_T_93 = {_ans_50_leadingZeros_T_49,_ans_50_leadingZeros_T_90,ans_50_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_50_leadingZeros_T_143 = _ans_50_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_144 = _ans_50_leadingZeros_T_93[46] ? 6'h2e : _ans_50_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_145 = _ans_50_leadingZeros_T_93[45] ? 6'h2d : _ans_50_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_146 = _ans_50_leadingZeros_T_93[44] ? 6'h2c : _ans_50_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_147 = _ans_50_leadingZeros_T_93[43] ? 6'h2b : _ans_50_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_148 = _ans_50_leadingZeros_T_93[42] ? 6'h2a : _ans_50_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_149 = _ans_50_leadingZeros_T_93[41] ? 6'h29 : _ans_50_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_150 = _ans_50_leadingZeros_T_93[40] ? 6'h28 : _ans_50_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_151 = _ans_50_leadingZeros_T_93[39] ? 6'h27 : _ans_50_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_152 = _ans_50_leadingZeros_T_93[38] ? 6'h26 : _ans_50_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_153 = _ans_50_leadingZeros_T_93[37] ? 6'h25 : _ans_50_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_154 = _ans_50_leadingZeros_T_93[36] ? 6'h24 : _ans_50_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_155 = _ans_50_leadingZeros_T_93[35] ? 6'h23 : _ans_50_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_156 = _ans_50_leadingZeros_T_93[34] ? 6'h22 : _ans_50_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_157 = _ans_50_leadingZeros_T_93[33] ? 6'h21 : _ans_50_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_158 = _ans_50_leadingZeros_T_93[32] ? 6'h20 : _ans_50_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_159 = _ans_50_leadingZeros_T_93[31] ? 6'h1f : _ans_50_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_160 = _ans_50_leadingZeros_T_93[30] ? 6'h1e : _ans_50_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_161 = _ans_50_leadingZeros_T_93[29] ? 6'h1d : _ans_50_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_162 = _ans_50_leadingZeros_T_93[28] ? 6'h1c : _ans_50_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_163 = _ans_50_leadingZeros_T_93[27] ? 6'h1b : _ans_50_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_164 = _ans_50_leadingZeros_T_93[26] ? 6'h1a : _ans_50_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_165 = _ans_50_leadingZeros_T_93[25] ? 6'h19 : _ans_50_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_166 = _ans_50_leadingZeros_T_93[24] ? 6'h18 : _ans_50_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_167 = _ans_50_leadingZeros_T_93[23] ? 6'h17 : _ans_50_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_168 = _ans_50_leadingZeros_T_93[22] ? 6'h16 : _ans_50_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_169 = _ans_50_leadingZeros_T_93[21] ? 6'h15 : _ans_50_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_170 = _ans_50_leadingZeros_T_93[20] ? 6'h14 : _ans_50_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_171 = _ans_50_leadingZeros_T_93[19] ? 6'h13 : _ans_50_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_172 = _ans_50_leadingZeros_T_93[18] ? 6'h12 : _ans_50_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_173 = _ans_50_leadingZeros_T_93[17] ? 6'h11 : _ans_50_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_174 = _ans_50_leadingZeros_T_93[16] ? 6'h10 : _ans_50_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_175 = _ans_50_leadingZeros_T_93[15] ? 6'hf : _ans_50_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_176 = _ans_50_leadingZeros_T_93[14] ? 6'he : _ans_50_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_177 = _ans_50_leadingZeros_T_93[13] ? 6'hd : _ans_50_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_178 = _ans_50_leadingZeros_T_93[12] ? 6'hc : _ans_50_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_179 = _ans_50_leadingZeros_T_93[11] ? 6'hb : _ans_50_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_180 = _ans_50_leadingZeros_T_93[10] ? 6'ha : _ans_50_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_181 = _ans_50_leadingZeros_T_93[9] ? 6'h9 : _ans_50_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_182 = _ans_50_leadingZeros_T_93[8] ? 6'h8 : _ans_50_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_183 = _ans_50_leadingZeros_T_93[7] ? 6'h7 : _ans_50_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_184 = _ans_50_leadingZeros_T_93[6] ? 6'h6 : _ans_50_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_185 = _ans_50_leadingZeros_T_93[5] ? 6'h5 : _ans_50_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_186 = _ans_50_leadingZeros_T_93[4] ? 6'h4 : _ans_50_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_187 = _ans_50_leadingZeros_T_93[3] ? 6'h3 : _ans_50_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_188 = _ans_50_leadingZeros_T_93[2] ? 6'h2 : _ans_50_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_leadingZeros_T_189 = _ans_50_leadingZeros_T_93[1] ? 6'h1 : _ans_50_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_50_leadingZeros = _ans_50_leadingZeros_T_93[0] ? 6'h0 : _ans_50_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_50_expRaw_T_1 = 6'h1f - ans_50_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_50_expRaw = ans_50_isZero ? 6'h0 : _ans_50_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_50_shiftAmt_T_2 = ans_50_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_50_shiftAmt = ans_50_expRaw > 6'h3 ? _ans_50_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_50_mantissaRaw_T = ans_50_absClipped >> ans_50_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_50_mantissaRaw = _ans_50_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_50_mantissa = ans_50_expRaw >= 6'h3 ? ans_50_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_50_expAdjusted = ans_50_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_50_exp_T_4 = ans_50_expAdjusted > 7'hf ? 4'hf : ans_50_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_50_exp = ans_50_isZero ? 4'h0 : _ans_50_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_50_fp8 = {ans_50_clippedX[31],ans_50_exp,ans_50_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_51 = {24'h0,linear_bias_51}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_51 = tempSum_51 + biasExtended_51; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_51_sign = sum32_51[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_51_absX_T = ~sum32_51; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_51_absX_T_2 = _ans_51_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_51_absX = ans_51_sign ? _ans_51_absX_T_2 : sum32_51; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_51_shiftedX_T_1 = _GEN_10432 - ans_51_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_51_shiftedX_T_3 = ans_51_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_51_shiftedX = ans_51_sign ? _ans_51_shiftedX_T_1 : _ans_51_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_51_scaledX_T_1 = ans_51_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_51_scaledX = _ans_51_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_51_clippedX_T_2 = ans_51_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_51_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_51_clippedX = ans_51_scaledX > 49'h1c0 ? 49'h1c0 : _ans_51_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_51_absClipped_T_1 = ~ans_51_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_51_absClipped_T_3 = _ans_51_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_51_absClipped = ans_51_clippedX[31] ? _ans_51_absClipped_T_3 : ans_51_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_51_isZero = ans_51_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_10995 = {{16'd0}, ans_51_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_4 = _GEN_10995 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_6 = {ans_51_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_8 = _ans_51_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_9 = _ans_51_leadingZeros_T_4 | _ans_51_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10996 = {{8'd0}, _ans_51_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_14 = _GEN_10996 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_16 = {_ans_51_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_18 = _ans_51_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_19 = _ans_51_leadingZeros_T_14 | _ans_51_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10997 = {{4'd0}, _ans_51_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_24 = _GEN_10997 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_26 = {_ans_51_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_28 = _ans_51_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_29 = _ans_51_leadingZeros_T_24 | _ans_51_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10998 = {{2'd0}, _ans_51_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_34 = _GEN_10998 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_36 = {_ans_51_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_38 = _ans_51_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_39 = _ans_51_leadingZeros_T_34 | _ans_51_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_10999 = {{1'd0}, _ans_51_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_44 = _GEN_10999 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_46 = {_ans_51_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_48 = _ans_51_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_51_leadingZeros_T_49 = _ans_51_leadingZeros_T_44 | _ans_51_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11000 = {{8'd0}, ans_51_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_55 = _GEN_11000 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_57 = {ans_51_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_59 = _ans_51_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_60 = _ans_51_leadingZeros_T_55 | _ans_51_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11001 = {{4'd0}, _ans_51_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_65 = _GEN_11001 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_67 = {_ans_51_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_69 = _ans_51_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_70 = _ans_51_leadingZeros_T_65 | _ans_51_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11002 = {{2'd0}, _ans_51_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_75 = _GEN_11002 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_77 = {_ans_51_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_79 = _ans_51_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_80 = _ans_51_leadingZeros_T_75 | _ans_51_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11003 = {{1'd0}, _ans_51_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_85 = _GEN_11003 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_87 = {_ans_51_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_89 = _ans_51_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_51_leadingZeros_T_90 = _ans_51_leadingZeros_T_85 | _ans_51_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_51_leadingZeros_T_93 = {_ans_51_leadingZeros_T_49,_ans_51_leadingZeros_T_90,ans_51_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_51_leadingZeros_T_143 = _ans_51_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_144 = _ans_51_leadingZeros_T_93[46] ? 6'h2e : _ans_51_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_145 = _ans_51_leadingZeros_T_93[45] ? 6'h2d : _ans_51_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_146 = _ans_51_leadingZeros_T_93[44] ? 6'h2c : _ans_51_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_147 = _ans_51_leadingZeros_T_93[43] ? 6'h2b : _ans_51_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_148 = _ans_51_leadingZeros_T_93[42] ? 6'h2a : _ans_51_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_149 = _ans_51_leadingZeros_T_93[41] ? 6'h29 : _ans_51_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_150 = _ans_51_leadingZeros_T_93[40] ? 6'h28 : _ans_51_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_151 = _ans_51_leadingZeros_T_93[39] ? 6'h27 : _ans_51_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_152 = _ans_51_leadingZeros_T_93[38] ? 6'h26 : _ans_51_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_153 = _ans_51_leadingZeros_T_93[37] ? 6'h25 : _ans_51_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_154 = _ans_51_leadingZeros_T_93[36] ? 6'h24 : _ans_51_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_155 = _ans_51_leadingZeros_T_93[35] ? 6'h23 : _ans_51_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_156 = _ans_51_leadingZeros_T_93[34] ? 6'h22 : _ans_51_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_157 = _ans_51_leadingZeros_T_93[33] ? 6'h21 : _ans_51_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_158 = _ans_51_leadingZeros_T_93[32] ? 6'h20 : _ans_51_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_159 = _ans_51_leadingZeros_T_93[31] ? 6'h1f : _ans_51_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_160 = _ans_51_leadingZeros_T_93[30] ? 6'h1e : _ans_51_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_161 = _ans_51_leadingZeros_T_93[29] ? 6'h1d : _ans_51_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_162 = _ans_51_leadingZeros_T_93[28] ? 6'h1c : _ans_51_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_163 = _ans_51_leadingZeros_T_93[27] ? 6'h1b : _ans_51_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_164 = _ans_51_leadingZeros_T_93[26] ? 6'h1a : _ans_51_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_165 = _ans_51_leadingZeros_T_93[25] ? 6'h19 : _ans_51_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_166 = _ans_51_leadingZeros_T_93[24] ? 6'h18 : _ans_51_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_167 = _ans_51_leadingZeros_T_93[23] ? 6'h17 : _ans_51_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_168 = _ans_51_leadingZeros_T_93[22] ? 6'h16 : _ans_51_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_169 = _ans_51_leadingZeros_T_93[21] ? 6'h15 : _ans_51_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_170 = _ans_51_leadingZeros_T_93[20] ? 6'h14 : _ans_51_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_171 = _ans_51_leadingZeros_T_93[19] ? 6'h13 : _ans_51_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_172 = _ans_51_leadingZeros_T_93[18] ? 6'h12 : _ans_51_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_173 = _ans_51_leadingZeros_T_93[17] ? 6'h11 : _ans_51_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_174 = _ans_51_leadingZeros_T_93[16] ? 6'h10 : _ans_51_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_175 = _ans_51_leadingZeros_T_93[15] ? 6'hf : _ans_51_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_176 = _ans_51_leadingZeros_T_93[14] ? 6'he : _ans_51_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_177 = _ans_51_leadingZeros_T_93[13] ? 6'hd : _ans_51_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_178 = _ans_51_leadingZeros_T_93[12] ? 6'hc : _ans_51_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_179 = _ans_51_leadingZeros_T_93[11] ? 6'hb : _ans_51_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_180 = _ans_51_leadingZeros_T_93[10] ? 6'ha : _ans_51_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_181 = _ans_51_leadingZeros_T_93[9] ? 6'h9 : _ans_51_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_182 = _ans_51_leadingZeros_T_93[8] ? 6'h8 : _ans_51_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_183 = _ans_51_leadingZeros_T_93[7] ? 6'h7 : _ans_51_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_184 = _ans_51_leadingZeros_T_93[6] ? 6'h6 : _ans_51_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_185 = _ans_51_leadingZeros_T_93[5] ? 6'h5 : _ans_51_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_186 = _ans_51_leadingZeros_T_93[4] ? 6'h4 : _ans_51_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_187 = _ans_51_leadingZeros_T_93[3] ? 6'h3 : _ans_51_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_188 = _ans_51_leadingZeros_T_93[2] ? 6'h2 : _ans_51_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_leadingZeros_T_189 = _ans_51_leadingZeros_T_93[1] ? 6'h1 : _ans_51_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_51_leadingZeros = _ans_51_leadingZeros_T_93[0] ? 6'h0 : _ans_51_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_51_expRaw_T_1 = 6'h1f - ans_51_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_51_expRaw = ans_51_isZero ? 6'h0 : _ans_51_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_51_shiftAmt_T_2 = ans_51_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_51_shiftAmt = ans_51_expRaw > 6'h3 ? _ans_51_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_51_mantissaRaw_T = ans_51_absClipped >> ans_51_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_51_mantissaRaw = _ans_51_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_51_mantissa = ans_51_expRaw >= 6'h3 ? ans_51_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_51_expAdjusted = ans_51_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_51_exp_T_4 = ans_51_expAdjusted > 7'hf ? 4'hf : ans_51_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_51_exp = ans_51_isZero ? 4'h0 : _ans_51_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_51_fp8 = {ans_51_clippedX[31],ans_51_exp,ans_51_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_52 = {24'h0,linear_bias_52}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_52 = tempSum_52 + biasExtended_52; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_52_sign = sum32_52[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_52_absX_T = ~sum32_52; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_52_absX_T_2 = _ans_52_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_52_absX = ans_52_sign ? _ans_52_absX_T_2 : sum32_52; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_52_shiftedX_T_1 = _GEN_10432 - ans_52_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_52_shiftedX_T_3 = ans_52_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_52_shiftedX = ans_52_sign ? _ans_52_shiftedX_T_1 : _ans_52_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_52_scaledX_T_1 = ans_52_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_52_scaledX = _ans_52_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_52_clippedX_T_2 = ans_52_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_52_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_52_clippedX = ans_52_scaledX > 49'h1c0 ? 49'h1c0 : _ans_52_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_52_absClipped_T_1 = ~ans_52_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_52_absClipped_T_3 = _ans_52_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_52_absClipped = ans_52_clippedX[31] ? _ans_52_absClipped_T_3 : ans_52_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_52_isZero = ans_52_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11006 = {{16'd0}, ans_52_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_4 = _GEN_11006 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_6 = {ans_52_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_8 = _ans_52_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_9 = _ans_52_leadingZeros_T_4 | _ans_52_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11007 = {{8'd0}, _ans_52_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_14 = _GEN_11007 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_16 = {_ans_52_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_18 = _ans_52_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_19 = _ans_52_leadingZeros_T_14 | _ans_52_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11008 = {{4'd0}, _ans_52_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_24 = _GEN_11008 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_26 = {_ans_52_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_28 = _ans_52_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_29 = _ans_52_leadingZeros_T_24 | _ans_52_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11009 = {{2'd0}, _ans_52_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_34 = _GEN_11009 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_36 = {_ans_52_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_38 = _ans_52_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_39 = _ans_52_leadingZeros_T_34 | _ans_52_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11010 = {{1'd0}, _ans_52_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_44 = _GEN_11010 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_46 = {_ans_52_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_48 = _ans_52_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_52_leadingZeros_T_49 = _ans_52_leadingZeros_T_44 | _ans_52_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11011 = {{8'd0}, ans_52_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_55 = _GEN_11011 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_57 = {ans_52_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_59 = _ans_52_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_60 = _ans_52_leadingZeros_T_55 | _ans_52_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11012 = {{4'd0}, _ans_52_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_65 = _GEN_11012 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_67 = {_ans_52_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_69 = _ans_52_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_70 = _ans_52_leadingZeros_T_65 | _ans_52_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11013 = {{2'd0}, _ans_52_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_75 = _GEN_11013 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_77 = {_ans_52_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_79 = _ans_52_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_80 = _ans_52_leadingZeros_T_75 | _ans_52_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11014 = {{1'd0}, _ans_52_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_85 = _GEN_11014 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_87 = {_ans_52_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_89 = _ans_52_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_52_leadingZeros_T_90 = _ans_52_leadingZeros_T_85 | _ans_52_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_52_leadingZeros_T_93 = {_ans_52_leadingZeros_T_49,_ans_52_leadingZeros_T_90,ans_52_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_52_leadingZeros_T_143 = _ans_52_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_144 = _ans_52_leadingZeros_T_93[46] ? 6'h2e : _ans_52_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_145 = _ans_52_leadingZeros_T_93[45] ? 6'h2d : _ans_52_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_146 = _ans_52_leadingZeros_T_93[44] ? 6'h2c : _ans_52_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_147 = _ans_52_leadingZeros_T_93[43] ? 6'h2b : _ans_52_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_148 = _ans_52_leadingZeros_T_93[42] ? 6'h2a : _ans_52_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_149 = _ans_52_leadingZeros_T_93[41] ? 6'h29 : _ans_52_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_150 = _ans_52_leadingZeros_T_93[40] ? 6'h28 : _ans_52_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_151 = _ans_52_leadingZeros_T_93[39] ? 6'h27 : _ans_52_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_152 = _ans_52_leadingZeros_T_93[38] ? 6'h26 : _ans_52_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_153 = _ans_52_leadingZeros_T_93[37] ? 6'h25 : _ans_52_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_154 = _ans_52_leadingZeros_T_93[36] ? 6'h24 : _ans_52_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_155 = _ans_52_leadingZeros_T_93[35] ? 6'h23 : _ans_52_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_156 = _ans_52_leadingZeros_T_93[34] ? 6'h22 : _ans_52_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_157 = _ans_52_leadingZeros_T_93[33] ? 6'h21 : _ans_52_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_158 = _ans_52_leadingZeros_T_93[32] ? 6'h20 : _ans_52_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_159 = _ans_52_leadingZeros_T_93[31] ? 6'h1f : _ans_52_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_160 = _ans_52_leadingZeros_T_93[30] ? 6'h1e : _ans_52_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_161 = _ans_52_leadingZeros_T_93[29] ? 6'h1d : _ans_52_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_162 = _ans_52_leadingZeros_T_93[28] ? 6'h1c : _ans_52_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_163 = _ans_52_leadingZeros_T_93[27] ? 6'h1b : _ans_52_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_164 = _ans_52_leadingZeros_T_93[26] ? 6'h1a : _ans_52_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_165 = _ans_52_leadingZeros_T_93[25] ? 6'h19 : _ans_52_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_166 = _ans_52_leadingZeros_T_93[24] ? 6'h18 : _ans_52_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_167 = _ans_52_leadingZeros_T_93[23] ? 6'h17 : _ans_52_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_168 = _ans_52_leadingZeros_T_93[22] ? 6'h16 : _ans_52_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_169 = _ans_52_leadingZeros_T_93[21] ? 6'h15 : _ans_52_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_170 = _ans_52_leadingZeros_T_93[20] ? 6'h14 : _ans_52_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_171 = _ans_52_leadingZeros_T_93[19] ? 6'h13 : _ans_52_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_172 = _ans_52_leadingZeros_T_93[18] ? 6'h12 : _ans_52_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_173 = _ans_52_leadingZeros_T_93[17] ? 6'h11 : _ans_52_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_174 = _ans_52_leadingZeros_T_93[16] ? 6'h10 : _ans_52_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_175 = _ans_52_leadingZeros_T_93[15] ? 6'hf : _ans_52_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_176 = _ans_52_leadingZeros_T_93[14] ? 6'he : _ans_52_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_177 = _ans_52_leadingZeros_T_93[13] ? 6'hd : _ans_52_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_178 = _ans_52_leadingZeros_T_93[12] ? 6'hc : _ans_52_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_179 = _ans_52_leadingZeros_T_93[11] ? 6'hb : _ans_52_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_180 = _ans_52_leadingZeros_T_93[10] ? 6'ha : _ans_52_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_181 = _ans_52_leadingZeros_T_93[9] ? 6'h9 : _ans_52_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_182 = _ans_52_leadingZeros_T_93[8] ? 6'h8 : _ans_52_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_183 = _ans_52_leadingZeros_T_93[7] ? 6'h7 : _ans_52_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_184 = _ans_52_leadingZeros_T_93[6] ? 6'h6 : _ans_52_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_185 = _ans_52_leadingZeros_T_93[5] ? 6'h5 : _ans_52_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_186 = _ans_52_leadingZeros_T_93[4] ? 6'h4 : _ans_52_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_187 = _ans_52_leadingZeros_T_93[3] ? 6'h3 : _ans_52_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_188 = _ans_52_leadingZeros_T_93[2] ? 6'h2 : _ans_52_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_leadingZeros_T_189 = _ans_52_leadingZeros_T_93[1] ? 6'h1 : _ans_52_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_52_leadingZeros = _ans_52_leadingZeros_T_93[0] ? 6'h0 : _ans_52_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_52_expRaw_T_1 = 6'h1f - ans_52_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_52_expRaw = ans_52_isZero ? 6'h0 : _ans_52_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_52_shiftAmt_T_2 = ans_52_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_52_shiftAmt = ans_52_expRaw > 6'h3 ? _ans_52_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_52_mantissaRaw_T = ans_52_absClipped >> ans_52_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_52_mantissaRaw = _ans_52_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_52_mantissa = ans_52_expRaw >= 6'h3 ? ans_52_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_52_expAdjusted = ans_52_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_52_exp_T_4 = ans_52_expAdjusted > 7'hf ? 4'hf : ans_52_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_52_exp = ans_52_isZero ? 4'h0 : _ans_52_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_52_fp8 = {ans_52_clippedX[31],ans_52_exp,ans_52_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_53 = {24'h0,linear_bias_53}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_53 = tempSum_53 + biasExtended_53; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_53_sign = sum32_53[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_53_absX_T = ~sum32_53; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_53_absX_T_2 = _ans_53_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_53_absX = ans_53_sign ? _ans_53_absX_T_2 : sum32_53; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_53_shiftedX_T_1 = _GEN_10432 - ans_53_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_53_shiftedX_T_3 = ans_53_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_53_shiftedX = ans_53_sign ? _ans_53_shiftedX_T_1 : _ans_53_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_53_scaledX_T_1 = ans_53_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_53_scaledX = _ans_53_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_53_clippedX_T_2 = ans_53_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_53_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_53_clippedX = ans_53_scaledX > 49'h1c0 ? 49'h1c0 : _ans_53_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_53_absClipped_T_1 = ~ans_53_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_53_absClipped_T_3 = _ans_53_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_53_absClipped = ans_53_clippedX[31] ? _ans_53_absClipped_T_3 : ans_53_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_53_isZero = ans_53_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11017 = {{16'd0}, ans_53_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_4 = _GEN_11017 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_6 = {ans_53_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_8 = _ans_53_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_9 = _ans_53_leadingZeros_T_4 | _ans_53_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11018 = {{8'd0}, _ans_53_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_14 = _GEN_11018 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_16 = {_ans_53_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_18 = _ans_53_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_19 = _ans_53_leadingZeros_T_14 | _ans_53_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11019 = {{4'd0}, _ans_53_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_24 = _GEN_11019 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_26 = {_ans_53_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_28 = _ans_53_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_29 = _ans_53_leadingZeros_T_24 | _ans_53_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11020 = {{2'd0}, _ans_53_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_34 = _GEN_11020 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_36 = {_ans_53_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_38 = _ans_53_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_39 = _ans_53_leadingZeros_T_34 | _ans_53_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11021 = {{1'd0}, _ans_53_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_44 = _GEN_11021 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_46 = {_ans_53_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_48 = _ans_53_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_53_leadingZeros_T_49 = _ans_53_leadingZeros_T_44 | _ans_53_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11022 = {{8'd0}, ans_53_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_55 = _GEN_11022 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_57 = {ans_53_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_59 = _ans_53_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_60 = _ans_53_leadingZeros_T_55 | _ans_53_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11023 = {{4'd0}, _ans_53_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_65 = _GEN_11023 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_67 = {_ans_53_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_69 = _ans_53_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_70 = _ans_53_leadingZeros_T_65 | _ans_53_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11024 = {{2'd0}, _ans_53_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_75 = _GEN_11024 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_77 = {_ans_53_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_79 = _ans_53_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_80 = _ans_53_leadingZeros_T_75 | _ans_53_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11025 = {{1'd0}, _ans_53_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_85 = _GEN_11025 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_87 = {_ans_53_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_89 = _ans_53_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_53_leadingZeros_T_90 = _ans_53_leadingZeros_T_85 | _ans_53_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_53_leadingZeros_T_93 = {_ans_53_leadingZeros_T_49,_ans_53_leadingZeros_T_90,ans_53_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_53_leadingZeros_T_143 = _ans_53_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_144 = _ans_53_leadingZeros_T_93[46] ? 6'h2e : _ans_53_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_145 = _ans_53_leadingZeros_T_93[45] ? 6'h2d : _ans_53_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_146 = _ans_53_leadingZeros_T_93[44] ? 6'h2c : _ans_53_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_147 = _ans_53_leadingZeros_T_93[43] ? 6'h2b : _ans_53_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_148 = _ans_53_leadingZeros_T_93[42] ? 6'h2a : _ans_53_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_149 = _ans_53_leadingZeros_T_93[41] ? 6'h29 : _ans_53_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_150 = _ans_53_leadingZeros_T_93[40] ? 6'h28 : _ans_53_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_151 = _ans_53_leadingZeros_T_93[39] ? 6'h27 : _ans_53_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_152 = _ans_53_leadingZeros_T_93[38] ? 6'h26 : _ans_53_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_153 = _ans_53_leadingZeros_T_93[37] ? 6'h25 : _ans_53_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_154 = _ans_53_leadingZeros_T_93[36] ? 6'h24 : _ans_53_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_155 = _ans_53_leadingZeros_T_93[35] ? 6'h23 : _ans_53_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_156 = _ans_53_leadingZeros_T_93[34] ? 6'h22 : _ans_53_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_157 = _ans_53_leadingZeros_T_93[33] ? 6'h21 : _ans_53_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_158 = _ans_53_leadingZeros_T_93[32] ? 6'h20 : _ans_53_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_159 = _ans_53_leadingZeros_T_93[31] ? 6'h1f : _ans_53_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_160 = _ans_53_leadingZeros_T_93[30] ? 6'h1e : _ans_53_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_161 = _ans_53_leadingZeros_T_93[29] ? 6'h1d : _ans_53_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_162 = _ans_53_leadingZeros_T_93[28] ? 6'h1c : _ans_53_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_163 = _ans_53_leadingZeros_T_93[27] ? 6'h1b : _ans_53_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_164 = _ans_53_leadingZeros_T_93[26] ? 6'h1a : _ans_53_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_165 = _ans_53_leadingZeros_T_93[25] ? 6'h19 : _ans_53_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_166 = _ans_53_leadingZeros_T_93[24] ? 6'h18 : _ans_53_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_167 = _ans_53_leadingZeros_T_93[23] ? 6'h17 : _ans_53_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_168 = _ans_53_leadingZeros_T_93[22] ? 6'h16 : _ans_53_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_169 = _ans_53_leadingZeros_T_93[21] ? 6'h15 : _ans_53_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_170 = _ans_53_leadingZeros_T_93[20] ? 6'h14 : _ans_53_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_171 = _ans_53_leadingZeros_T_93[19] ? 6'h13 : _ans_53_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_172 = _ans_53_leadingZeros_T_93[18] ? 6'h12 : _ans_53_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_173 = _ans_53_leadingZeros_T_93[17] ? 6'h11 : _ans_53_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_174 = _ans_53_leadingZeros_T_93[16] ? 6'h10 : _ans_53_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_175 = _ans_53_leadingZeros_T_93[15] ? 6'hf : _ans_53_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_176 = _ans_53_leadingZeros_T_93[14] ? 6'he : _ans_53_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_177 = _ans_53_leadingZeros_T_93[13] ? 6'hd : _ans_53_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_178 = _ans_53_leadingZeros_T_93[12] ? 6'hc : _ans_53_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_179 = _ans_53_leadingZeros_T_93[11] ? 6'hb : _ans_53_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_180 = _ans_53_leadingZeros_T_93[10] ? 6'ha : _ans_53_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_181 = _ans_53_leadingZeros_T_93[9] ? 6'h9 : _ans_53_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_182 = _ans_53_leadingZeros_T_93[8] ? 6'h8 : _ans_53_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_183 = _ans_53_leadingZeros_T_93[7] ? 6'h7 : _ans_53_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_184 = _ans_53_leadingZeros_T_93[6] ? 6'h6 : _ans_53_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_185 = _ans_53_leadingZeros_T_93[5] ? 6'h5 : _ans_53_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_186 = _ans_53_leadingZeros_T_93[4] ? 6'h4 : _ans_53_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_187 = _ans_53_leadingZeros_T_93[3] ? 6'h3 : _ans_53_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_188 = _ans_53_leadingZeros_T_93[2] ? 6'h2 : _ans_53_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_leadingZeros_T_189 = _ans_53_leadingZeros_T_93[1] ? 6'h1 : _ans_53_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_53_leadingZeros = _ans_53_leadingZeros_T_93[0] ? 6'h0 : _ans_53_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_53_expRaw_T_1 = 6'h1f - ans_53_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_53_expRaw = ans_53_isZero ? 6'h0 : _ans_53_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_53_shiftAmt_T_2 = ans_53_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_53_shiftAmt = ans_53_expRaw > 6'h3 ? _ans_53_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_53_mantissaRaw_T = ans_53_absClipped >> ans_53_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_53_mantissaRaw = _ans_53_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_53_mantissa = ans_53_expRaw >= 6'h3 ? ans_53_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_53_expAdjusted = ans_53_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_53_exp_T_4 = ans_53_expAdjusted > 7'hf ? 4'hf : ans_53_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_53_exp = ans_53_isZero ? 4'h0 : _ans_53_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_53_fp8 = {ans_53_clippedX[31],ans_53_exp,ans_53_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_54 = {24'h0,linear_bias_54}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_54 = tempSum_54 + biasExtended_54; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_54_sign = sum32_54[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_54_absX_T = ~sum32_54; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_54_absX_T_2 = _ans_54_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_54_absX = ans_54_sign ? _ans_54_absX_T_2 : sum32_54; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_54_shiftedX_T_1 = _GEN_10432 - ans_54_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_54_shiftedX_T_3 = ans_54_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_54_shiftedX = ans_54_sign ? _ans_54_shiftedX_T_1 : _ans_54_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_54_scaledX_T_1 = ans_54_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_54_scaledX = _ans_54_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_54_clippedX_T_2 = ans_54_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_54_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_54_clippedX = ans_54_scaledX > 49'h1c0 ? 49'h1c0 : _ans_54_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_54_absClipped_T_1 = ~ans_54_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_54_absClipped_T_3 = _ans_54_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_54_absClipped = ans_54_clippedX[31] ? _ans_54_absClipped_T_3 : ans_54_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_54_isZero = ans_54_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11028 = {{16'd0}, ans_54_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_4 = _GEN_11028 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_6 = {ans_54_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_8 = _ans_54_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_9 = _ans_54_leadingZeros_T_4 | _ans_54_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11029 = {{8'd0}, _ans_54_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_14 = _GEN_11029 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_16 = {_ans_54_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_18 = _ans_54_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_19 = _ans_54_leadingZeros_T_14 | _ans_54_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11030 = {{4'd0}, _ans_54_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_24 = _GEN_11030 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_26 = {_ans_54_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_28 = _ans_54_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_29 = _ans_54_leadingZeros_T_24 | _ans_54_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11031 = {{2'd0}, _ans_54_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_34 = _GEN_11031 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_36 = {_ans_54_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_38 = _ans_54_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_39 = _ans_54_leadingZeros_T_34 | _ans_54_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11032 = {{1'd0}, _ans_54_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_44 = _GEN_11032 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_46 = {_ans_54_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_48 = _ans_54_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_54_leadingZeros_T_49 = _ans_54_leadingZeros_T_44 | _ans_54_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11033 = {{8'd0}, ans_54_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_55 = _GEN_11033 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_57 = {ans_54_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_59 = _ans_54_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_60 = _ans_54_leadingZeros_T_55 | _ans_54_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11034 = {{4'd0}, _ans_54_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_65 = _GEN_11034 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_67 = {_ans_54_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_69 = _ans_54_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_70 = _ans_54_leadingZeros_T_65 | _ans_54_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11035 = {{2'd0}, _ans_54_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_75 = _GEN_11035 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_77 = {_ans_54_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_79 = _ans_54_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_80 = _ans_54_leadingZeros_T_75 | _ans_54_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11036 = {{1'd0}, _ans_54_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_85 = _GEN_11036 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_87 = {_ans_54_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_89 = _ans_54_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_54_leadingZeros_T_90 = _ans_54_leadingZeros_T_85 | _ans_54_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_54_leadingZeros_T_93 = {_ans_54_leadingZeros_T_49,_ans_54_leadingZeros_T_90,ans_54_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_54_leadingZeros_T_143 = _ans_54_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_144 = _ans_54_leadingZeros_T_93[46] ? 6'h2e : _ans_54_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_145 = _ans_54_leadingZeros_T_93[45] ? 6'h2d : _ans_54_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_146 = _ans_54_leadingZeros_T_93[44] ? 6'h2c : _ans_54_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_147 = _ans_54_leadingZeros_T_93[43] ? 6'h2b : _ans_54_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_148 = _ans_54_leadingZeros_T_93[42] ? 6'h2a : _ans_54_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_149 = _ans_54_leadingZeros_T_93[41] ? 6'h29 : _ans_54_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_150 = _ans_54_leadingZeros_T_93[40] ? 6'h28 : _ans_54_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_151 = _ans_54_leadingZeros_T_93[39] ? 6'h27 : _ans_54_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_152 = _ans_54_leadingZeros_T_93[38] ? 6'h26 : _ans_54_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_153 = _ans_54_leadingZeros_T_93[37] ? 6'h25 : _ans_54_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_154 = _ans_54_leadingZeros_T_93[36] ? 6'h24 : _ans_54_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_155 = _ans_54_leadingZeros_T_93[35] ? 6'h23 : _ans_54_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_156 = _ans_54_leadingZeros_T_93[34] ? 6'h22 : _ans_54_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_157 = _ans_54_leadingZeros_T_93[33] ? 6'h21 : _ans_54_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_158 = _ans_54_leadingZeros_T_93[32] ? 6'h20 : _ans_54_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_159 = _ans_54_leadingZeros_T_93[31] ? 6'h1f : _ans_54_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_160 = _ans_54_leadingZeros_T_93[30] ? 6'h1e : _ans_54_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_161 = _ans_54_leadingZeros_T_93[29] ? 6'h1d : _ans_54_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_162 = _ans_54_leadingZeros_T_93[28] ? 6'h1c : _ans_54_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_163 = _ans_54_leadingZeros_T_93[27] ? 6'h1b : _ans_54_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_164 = _ans_54_leadingZeros_T_93[26] ? 6'h1a : _ans_54_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_165 = _ans_54_leadingZeros_T_93[25] ? 6'h19 : _ans_54_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_166 = _ans_54_leadingZeros_T_93[24] ? 6'h18 : _ans_54_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_167 = _ans_54_leadingZeros_T_93[23] ? 6'h17 : _ans_54_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_168 = _ans_54_leadingZeros_T_93[22] ? 6'h16 : _ans_54_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_169 = _ans_54_leadingZeros_T_93[21] ? 6'h15 : _ans_54_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_170 = _ans_54_leadingZeros_T_93[20] ? 6'h14 : _ans_54_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_171 = _ans_54_leadingZeros_T_93[19] ? 6'h13 : _ans_54_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_172 = _ans_54_leadingZeros_T_93[18] ? 6'h12 : _ans_54_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_173 = _ans_54_leadingZeros_T_93[17] ? 6'h11 : _ans_54_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_174 = _ans_54_leadingZeros_T_93[16] ? 6'h10 : _ans_54_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_175 = _ans_54_leadingZeros_T_93[15] ? 6'hf : _ans_54_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_176 = _ans_54_leadingZeros_T_93[14] ? 6'he : _ans_54_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_177 = _ans_54_leadingZeros_T_93[13] ? 6'hd : _ans_54_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_178 = _ans_54_leadingZeros_T_93[12] ? 6'hc : _ans_54_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_179 = _ans_54_leadingZeros_T_93[11] ? 6'hb : _ans_54_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_180 = _ans_54_leadingZeros_T_93[10] ? 6'ha : _ans_54_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_181 = _ans_54_leadingZeros_T_93[9] ? 6'h9 : _ans_54_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_182 = _ans_54_leadingZeros_T_93[8] ? 6'h8 : _ans_54_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_183 = _ans_54_leadingZeros_T_93[7] ? 6'h7 : _ans_54_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_184 = _ans_54_leadingZeros_T_93[6] ? 6'h6 : _ans_54_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_185 = _ans_54_leadingZeros_T_93[5] ? 6'h5 : _ans_54_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_186 = _ans_54_leadingZeros_T_93[4] ? 6'h4 : _ans_54_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_187 = _ans_54_leadingZeros_T_93[3] ? 6'h3 : _ans_54_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_188 = _ans_54_leadingZeros_T_93[2] ? 6'h2 : _ans_54_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_leadingZeros_T_189 = _ans_54_leadingZeros_T_93[1] ? 6'h1 : _ans_54_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_54_leadingZeros = _ans_54_leadingZeros_T_93[0] ? 6'h0 : _ans_54_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_54_expRaw_T_1 = 6'h1f - ans_54_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_54_expRaw = ans_54_isZero ? 6'h0 : _ans_54_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_54_shiftAmt_T_2 = ans_54_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_54_shiftAmt = ans_54_expRaw > 6'h3 ? _ans_54_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_54_mantissaRaw_T = ans_54_absClipped >> ans_54_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_54_mantissaRaw = _ans_54_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_54_mantissa = ans_54_expRaw >= 6'h3 ? ans_54_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_54_expAdjusted = ans_54_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_54_exp_T_4 = ans_54_expAdjusted > 7'hf ? 4'hf : ans_54_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_54_exp = ans_54_isZero ? 4'h0 : _ans_54_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_54_fp8 = {ans_54_clippedX[31],ans_54_exp,ans_54_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_55 = {24'h0,linear_bias_55}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_55 = tempSum_55 + biasExtended_55; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_55_sign = sum32_55[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_55_absX_T = ~sum32_55; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_55_absX_T_2 = _ans_55_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_55_absX = ans_55_sign ? _ans_55_absX_T_2 : sum32_55; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_55_shiftedX_T_1 = _GEN_10432 - ans_55_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_55_shiftedX_T_3 = ans_55_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_55_shiftedX = ans_55_sign ? _ans_55_shiftedX_T_1 : _ans_55_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_55_scaledX_T_1 = ans_55_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_55_scaledX = _ans_55_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_55_clippedX_T_2 = ans_55_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_55_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_55_clippedX = ans_55_scaledX > 49'h1c0 ? 49'h1c0 : _ans_55_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_55_absClipped_T_1 = ~ans_55_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_55_absClipped_T_3 = _ans_55_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_55_absClipped = ans_55_clippedX[31] ? _ans_55_absClipped_T_3 : ans_55_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_55_isZero = ans_55_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11039 = {{16'd0}, ans_55_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_4 = _GEN_11039 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_6 = {ans_55_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_8 = _ans_55_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_9 = _ans_55_leadingZeros_T_4 | _ans_55_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11040 = {{8'd0}, _ans_55_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_14 = _GEN_11040 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_16 = {_ans_55_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_18 = _ans_55_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_19 = _ans_55_leadingZeros_T_14 | _ans_55_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11041 = {{4'd0}, _ans_55_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_24 = _GEN_11041 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_26 = {_ans_55_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_28 = _ans_55_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_29 = _ans_55_leadingZeros_T_24 | _ans_55_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11042 = {{2'd0}, _ans_55_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_34 = _GEN_11042 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_36 = {_ans_55_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_38 = _ans_55_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_39 = _ans_55_leadingZeros_T_34 | _ans_55_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11043 = {{1'd0}, _ans_55_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_44 = _GEN_11043 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_46 = {_ans_55_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_48 = _ans_55_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_55_leadingZeros_T_49 = _ans_55_leadingZeros_T_44 | _ans_55_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11044 = {{8'd0}, ans_55_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_55 = _GEN_11044 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_57 = {ans_55_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_59 = _ans_55_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_60 = _ans_55_leadingZeros_T_55 | _ans_55_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11045 = {{4'd0}, _ans_55_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_65 = _GEN_11045 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_67 = {_ans_55_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_69 = _ans_55_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_70 = _ans_55_leadingZeros_T_65 | _ans_55_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11046 = {{2'd0}, _ans_55_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_75 = _GEN_11046 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_77 = {_ans_55_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_79 = _ans_55_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_80 = _ans_55_leadingZeros_T_75 | _ans_55_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11047 = {{1'd0}, _ans_55_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_85 = _GEN_11047 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_87 = {_ans_55_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_89 = _ans_55_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_55_leadingZeros_T_90 = _ans_55_leadingZeros_T_85 | _ans_55_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_55_leadingZeros_T_93 = {_ans_55_leadingZeros_T_49,_ans_55_leadingZeros_T_90,ans_55_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_55_leadingZeros_T_143 = _ans_55_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_144 = _ans_55_leadingZeros_T_93[46] ? 6'h2e : _ans_55_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_145 = _ans_55_leadingZeros_T_93[45] ? 6'h2d : _ans_55_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_146 = _ans_55_leadingZeros_T_93[44] ? 6'h2c : _ans_55_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_147 = _ans_55_leadingZeros_T_93[43] ? 6'h2b : _ans_55_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_148 = _ans_55_leadingZeros_T_93[42] ? 6'h2a : _ans_55_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_149 = _ans_55_leadingZeros_T_93[41] ? 6'h29 : _ans_55_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_150 = _ans_55_leadingZeros_T_93[40] ? 6'h28 : _ans_55_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_151 = _ans_55_leadingZeros_T_93[39] ? 6'h27 : _ans_55_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_152 = _ans_55_leadingZeros_T_93[38] ? 6'h26 : _ans_55_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_153 = _ans_55_leadingZeros_T_93[37] ? 6'h25 : _ans_55_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_154 = _ans_55_leadingZeros_T_93[36] ? 6'h24 : _ans_55_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_155 = _ans_55_leadingZeros_T_93[35] ? 6'h23 : _ans_55_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_156 = _ans_55_leadingZeros_T_93[34] ? 6'h22 : _ans_55_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_157 = _ans_55_leadingZeros_T_93[33] ? 6'h21 : _ans_55_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_158 = _ans_55_leadingZeros_T_93[32] ? 6'h20 : _ans_55_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_159 = _ans_55_leadingZeros_T_93[31] ? 6'h1f : _ans_55_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_160 = _ans_55_leadingZeros_T_93[30] ? 6'h1e : _ans_55_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_161 = _ans_55_leadingZeros_T_93[29] ? 6'h1d : _ans_55_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_162 = _ans_55_leadingZeros_T_93[28] ? 6'h1c : _ans_55_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_163 = _ans_55_leadingZeros_T_93[27] ? 6'h1b : _ans_55_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_164 = _ans_55_leadingZeros_T_93[26] ? 6'h1a : _ans_55_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_165 = _ans_55_leadingZeros_T_93[25] ? 6'h19 : _ans_55_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_166 = _ans_55_leadingZeros_T_93[24] ? 6'h18 : _ans_55_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_167 = _ans_55_leadingZeros_T_93[23] ? 6'h17 : _ans_55_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_168 = _ans_55_leadingZeros_T_93[22] ? 6'h16 : _ans_55_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_169 = _ans_55_leadingZeros_T_93[21] ? 6'h15 : _ans_55_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_170 = _ans_55_leadingZeros_T_93[20] ? 6'h14 : _ans_55_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_171 = _ans_55_leadingZeros_T_93[19] ? 6'h13 : _ans_55_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_172 = _ans_55_leadingZeros_T_93[18] ? 6'h12 : _ans_55_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_173 = _ans_55_leadingZeros_T_93[17] ? 6'h11 : _ans_55_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_174 = _ans_55_leadingZeros_T_93[16] ? 6'h10 : _ans_55_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_175 = _ans_55_leadingZeros_T_93[15] ? 6'hf : _ans_55_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_176 = _ans_55_leadingZeros_T_93[14] ? 6'he : _ans_55_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_177 = _ans_55_leadingZeros_T_93[13] ? 6'hd : _ans_55_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_178 = _ans_55_leadingZeros_T_93[12] ? 6'hc : _ans_55_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_179 = _ans_55_leadingZeros_T_93[11] ? 6'hb : _ans_55_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_180 = _ans_55_leadingZeros_T_93[10] ? 6'ha : _ans_55_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_181 = _ans_55_leadingZeros_T_93[9] ? 6'h9 : _ans_55_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_182 = _ans_55_leadingZeros_T_93[8] ? 6'h8 : _ans_55_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_183 = _ans_55_leadingZeros_T_93[7] ? 6'h7 : _ans_55_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_184 = _ans_55_leadingZeros_T_93[6] ? 6'h6 : _ans_55_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_185 = _ans_55_leadingZeros_T_93[5] ? 6'h5 : _ans_55_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_186 = _ans_55_leadingZeros_T_93[4] ? 6'h4 : _ans_55_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_187 = _ans_55_leadingZeros_T_93[3] ? 6'h3 : _ans_55_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_188 = _ans_55_leadingZeros_T_93[2] ? 6'h2 : _ans_55_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_leadingZeros_T_189 = _ans_55_leadingZeros_T_93[1] ? 6'h1 : _ans_55_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_55_leadingZeros = _ans_55_leadingZeros_T_93[0] ? 6'h0 : _ans_55_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_55_expRaw_T_1 = 6'h1f - ans_55_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_55_expRaw = ans_55_isZero ? 6'h0 : _ans_55_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_55_shiftAmt_T_2 = ans_55_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_55_shiftAmt = ans_55_expRaw > 6'h3 ? _ans_55_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_55_mantissaRaw_T = ans_55_absClipped >> ans_55_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_55_mantissaRaw = _ans_55_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_55_mantissa = ans_55_expRaw >= 6'h3 ? ans_55_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_55_expAdjusted = ans_55_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_55_exp_T_4 = ans_55_expAdjusted > 7'hf ? 4'hf : ans_55_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_55_exp = ans_55_isZero ? 4'h0 : _ans_55_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_55_fp8 = {ans_55_clippedX[31],ans_55_exp,ans_55_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_56 = {24'h0,linear_bias_56}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_56 = tempSum_56 + biasExtended_56; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_56_sign = sum32_56[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_56_absX_T = ~sum32_56; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_56_absX_T_2 = _ans_56_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_56_absX = ans_56_sign ? _ans_56_absX_T_2 : sum32_56; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_56_shiftedX_T_1 = _GEN_10432 - ans_56_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_56_shiftedX_T_3 = ans_56_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_56_shiftedX = ans_56_sign ? _ans_56_shiftedX_T_1 : _ans_56_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_56_scaledX_T_1 = ans_56_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_56_scaledX = _ans_56_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_56_clippedX_T_2 = ans_56_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_56_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_56_clippedX = ans_56_scaledX > 49'h1c0 ? 49'h1c0 : _ans_56_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_56_absClipped_T_1 = ~ans_56_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_56_absClipped_T_3 = _ans_56_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_56_absClipped = ans_56_clippedX[31] ? _ans_56_absClipped_T_3 : ans_56_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_56_isZero = ans_56_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11050 = {{16'd0}, ans_56_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_4 = _GEN_11050 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_6 = {ans_56_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_8 = _ans_56_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_9 = _ans_56_leadingZeros_T_4 | _ans_56_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11051 = {{8'd0}, _ans_56_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_14 = _GEN_11051 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_16 = {_ans_56_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_18 = _ans_56_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_19 = _ans_56_leadingZeros_T_14 | _ans_56_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11052 = {{4'd0}, _ans_56_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_24 = _GEN_11052 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_26 = {_ans_56_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_28 = _ans_56_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_29 = _ans_56_leadingZeros_T_24 | _ans_56_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11053 = {{2'd0}, _ans_56_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_34 = _GEN_11053 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_36 = {_ans_56_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_38 = _ans_56_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_39 = _ans_56_leadingZeros_T_34 | _ans_56_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11054 = {{1'd0}, _ans_56_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_44 = _GEN_11054 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_46 = {_ans_56_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_48 = _ans_56_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_56_leadingZeros_T_49 = _ans_56_leadingZeros_T_44 | _ans_56_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11055 = {{8'd0}, ans_56_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_55 = _GEN_11055 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_57 = {ans_56_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_59 = _ans_56_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_60 = _ans_56_leadingZeros_T_55 | _ans_56_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11056 = {{4'd0}, _ans_56_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_65 = _GEN_11056 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_67 = {_ans_56_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_69 = _ans_56_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_70 = _ans_56_leadingZeros_T_65 | _ans_56_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11057 = {{2'd0}, _ans_56_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_75 = _GEN_11057 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_77 = {_ans_56_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_79 = _ans_56_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_80 = _ans_56_leadingZeros_T_75 | _ans_56_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11058 = {{1'd0}, _ans_56_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_85 = _GEN_11058 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_87 = {_ans_56_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_89 = _ans_56_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_56_leadingZeros_T_90 = _ans_56_leadingZeros_T_85 | _ans_56_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_56_leadingZeros_T_93 = {_ans_56_leadingZeros_T_49,_ans_56_leadingZeros_T_90,ans_56_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_56_leadingZeros_T_143 = _ans_56_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_144 = _ans_56_leadingZeros_T_93[46] ? 6'h2e : _ans_56_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_145 = _ans_56_leadingZeros_T_93[45] ? 6'h2d : _ans_56_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_146 = _ans_56_leadingZeros_T_93[44] ? 6'h2c : _ans_56_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_147 = _ans_56_leadingZeros_T_93[43] ? 6'h2b : _ans_56_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_148 = _ans_56_leadingZeros_T_93[42] ? 6'h2a : _ans_56_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_149 = _ans_56_leadingZeros_T_93[41] ? 6'h29 : _ans_56_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_150 = _ans_56_leadingZeros_T_93[40] ? 6'h28 : _ans_56_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_151 = _ans_56_leadingZeros_T_93[39] ? 6'h27 : _ans_56_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_152 = _ans_56_leadingZeros_T_93[38] ? 6'h26 : _ans_56_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_153 = _ans_56_leadingZeros_T_93[37] ? 6'h25 : _ans_56_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_154 = _ans_56_leadingZeros_T_93[36] ? 6'h24 : _ans_56_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_155 = _ans_56_leadingZeros_T_93[35] ? 6'h23 : _ans_56_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_156 = _ans_56_leadingZeros_T_93[34] ? 6'h22 : _ans_56_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_157 = _ans_56_leadingZeros_T_93[33] ? 6'h21 : _ans_56_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_158 = _ans_56_leadingZeros_T_93[32] ? 6'h20 : _ans_56_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_159 = _ans_56_leadingZeros_T_93[31] ? 6'h1f : _ans_56_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_160 = _ans_56_leadingZeros_T_93[30] ? 6'h1e : _ans_56_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_161 = _ans_56_leadingZeros_T_93[29] ? 6'h1d : _ans_56_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_162 = _ans_56_leadingZeros_T_93[28] ? 6'h1c : _ans_56_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_163 = _ans_56_leadingZeros_T_93[27] ? 6'h1b : _ans_56_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_164 = _ans_56_leadingZeros_T_93[26] ? 6'h1a : _ans_56_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_165 = _ans_56_leadingZeros_T_93[25] ? 6'h19 : _ans_56_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_166 = _ans_56_leadingZeros_T_93[24] ? 6'h18 : _ans_56_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_167 = _ans_56_leadingZeros_T_93[23] ? 6'h17 : _ans_56_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_168 = _ans_56_leadingZeros_T_93[22] ? 6'h16 : _ans_56_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_169 = _ans_56_leadingZeros_T_93[21] ? 6'h15 : _ans_56_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_170 = _ans_56_leadingZeros_T_93[20] ? 6'h14 : _ans_56_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_171 = _ans_56_leadingZeros_T_93[19] ? 6'h13 : _ans_56_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_172 = _ans_56_leadingZeros_T_93[18] ? 6'h12 : _ans_56_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_173 = _ans_56_leadingZeros_T_93[17] ? 6'h11 : _ans_56_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_174 = _ans_56_leadingZeros_T_93[16] ? 6'h10 : _ans_56_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_175 = _ans_56_leadingZeros_T_93[15] ? 6'hf : _ans_56_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_176 = _ans_56_leadingZeros_T_93[14] ? 6'he : _ans_56_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_177 = _ans_56_leadingZeros_T_93[13] ? 6'hd : _ans_56_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_178 = _ans_56_leadingZeros_T_93[12] ? 6'hc : _ans_56_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_179 = _ans_56_leadingZeros_T_93[11] ? 6'hb : _ans_56_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_180 = _ans_56_leadingZeros_T_93[10] ? 6'ha : _ans_56_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_181 = _ans_56_leadingZeros_T_93[9] ? 6'h9 : _ans_56_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_182 = _ans_56_leadingZeros_T_93[8] ? 6'h8 : _ans_56_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_183 = _ans_56_leadingZeros_T_93[7] ? 6'h7 : _ans_56_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_184 = _ans_56_leadingZeros_T_93[6] ? 6'h6 : _ans_56_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_185 = _ans_56_leadingZeros_T_93[5] ? 6'h5 : _ans_56_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_186 = _ans_56_leadingZeros_T_93[4] ? 6'h4 : _ans_56_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_187 = _ans_56_leadingZeros_T_93[3] ? 6'h3 : _ans_56_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_188 = _ans_56_leadingZeros_T_93[2] ? 6'h2 : _ans_56_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_leadingZeros_T_189 = _ans_56_leadingZeros_T_93[1] ? 6'h1 : _ans_56_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_56_leadingZeros = _ans_56_leadingZeros_T_93[0] ? 6'h0 : _ans_56_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_56_expRaw_T_1 = 6'h1f - ans_56_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_56_expRaw = ans_56_isZero ? 6'h0 : _ans_56_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_56_shiftAmt_T_2 = ans_56_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_56_shiftAmt = ans_56_expRaw > 6'h3 ? _ans_56_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_56_mantissaRaw_T = ans_56_absClipped >> ans_56_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_56_mantissaRaw = _ans_56_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_56_mantissa = ans_56_expRaw >= 6'h3 ? ans_56_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_56_expAdjusted = ans_56_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_56_exp_T_4 = ans_56_expAdjusted > 7'hf ? 4'hf : ans_56_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_56_exp = ans_56_isZero ? 4'h0 : _ans_56_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_56_fp8 = {ans_56_clippedX[31],ans_56_exp,ans_56_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_57 = {24'h0,linear_bias_57}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_57 = tempSum_57 + biasExtended_57; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_57_sign = sum32_57[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_57_absX_T = ~sum32_57; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_57_absX_T_2 = _ans_57_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_57_absX = ans_57_sign ? _ans_57_absX_T_2 : sum32_57; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_57_shiftedX_T_1 = _GEN_10432 - ans_57_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_57_shiftedX_T_3 = ans_57_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_57_shiftedX = ans_57_sign ? _ans_57_shiftedX_T_1 : _ans_57_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_57_scaledX_T_1 = ans_57_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_57_scaledX = _ans_57_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_57_clippedX_T_2 = ans_57_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_57_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_57_clippedX = ans_57_scaledX > 49'h1c0 ? 49'h1c0 : _ans_57_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_57_absClipped_T_1 = ~ans_57_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_57_absClipped_T_3 = _ans_57_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_57_absClipped = ans_57_clippedX[31] ? _ans_57_absClipped_T_3 : ans_57_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_57_isZero = ans_57_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11061 = {{16'd0}, ans_57_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_4 = _GEN_11061 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_6 = {ans_57_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_8 = _ans_57_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_9 = _ans_57_leadingZeros_T_4 | _ans_57_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11062 = {{8'd0}, _ans_57_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_14 = _GEN_11062 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_16 = {_ans_57_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_18 = _ans_57_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_19 = _ans_57_leadingZeros_T_14 | _ans_57_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11063 = {{4'd0}, _ans_57_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_24 = _GEN_11063 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_26 = {_ans_57_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_28 = _ans_57_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_29 = _ans_57_leadingZeros_T_24 | _ans_57_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11064 = {{2'd0}, _ans_57_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_34 = _GEN_11064 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_36 = {_ans_57_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_38 = _ans_57_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_39 = _ans_57_leadingZeros_T_34 | _ans_57_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11065 = {{1'd0}, _ans_57_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_44 = _GEN_11065 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_46 = {_ans_57_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_48 = _ans_57_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_57_leadingZeros_T_49 = _ans_57_leadingZeros_T_44 | _ans_57_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11066 = {{8'd0}, ans_57_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_55 = _GEN_11066 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_57 = {ans_57_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_59 = _ans_57_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_60 = _ans_57_leadingZeros_T_55 | _ans_57_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11067 = {{4'd0}, _ans_57_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_65 = _GEN_11067 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_67 = {_ans_57_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_69 = _ans_57_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_70 = _ans_57_leadingZeros_T_65 | _ans_57_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11068 = {{2'd0}, _ans_57_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_75 = _GEN_11068 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_77 = {_ans_57_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_79 = _ans_57_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_80 = _ans_57_leadingZeros_T_75 | _ans_57_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11069 = {{1'd0}, _ans_57_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_85 = _GEN_11069 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_87 = {_ans_57_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_89 = _ans_57_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_57_leadingZeros_T_90 = _ans_57_leadingZeros_T_85 | _ans_57_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_57_leadingZeros_T_93 = {_ans_57_leadingZeros_T_49,_ans_57_leadingZeros_T_90,ans_57_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_57_leadingZeros_T_143 = _ans_57_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_144 = _ans_57_leadingZeros_T_93[46] ? 6'h2e : _ans_57_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_145 = _ans_57_leadingZeros_T_93[45] ? 6'h2d : _ans_57_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_146 = _ans_57_leadingZeros_T_93[44] ? 6'h2c : _ans_57_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_147 = _ans_57_leadingZeros_T_93[43] ? 6'h2b : _ans_57_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_148 = _ans_57_leadingZeros_T_93[42] ? 6'h2a : _ans_57_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_149 = _ans_57_leadingZeros_T_93[41] ? 6'h29 : _ans_57_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_150 = _ans_57_leadingZeros_T_93[40] ? 6'h28 : _ans_57_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_151 = _ans_57_leadingZeros_T_93[39] ? 6'h27 : _ans_57_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_152 = _ans_57_leadingZeros_T_93[38] ? 6'h26 : _ans_57_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_153 = _ans_57_leadingZeros_T_93[37] ? 6'h25 : _ans_57_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_154 = _ans_57_leadingZeros_T_93[36] ? 6'h24 : _ans_57_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_155 = _ans_57_leadingZeros_T_93[35] ? 6'h23 : _ans_57_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_156 = _ans_57_leadingZeros_T_93[34] ? 6'h22 : _ans_57_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_157 = _ans_57_leadingZeros_T_93[33] ? 6'h21 : _ans_57_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_158 = _ans_57_leadingZeros_T_93[32] ? 6'h20 : _ans_57_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_159 = _ans_57_leadingZeros_T_93[31] ? 6'h1f : _ans_57_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_160 = _ans_57_leadingZeros_T_93[30] ? 6'h1e : _ans_57_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_161 = _ans_57_leadingZeros_T_93[29] ? 6'h1d : _ans_57_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_162 = _ans_57_leadingZeros_T_93[28] ? 6'h1c : _ans_57_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_163 = _ans_57_leadingZeros_T_93[27] ? 6'h1b : _ans_57_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_164 = _ans_57_leadingZeros_T_93[26] ? 6'h1a : _ans_57_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_165 = _ans_57_leadingZeros_T_93[25] ? 6'h19 : _ans_57_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_166 = _ans_57_leadingZeros_T_93[24] ? 6'h18 : _ans_57_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_167 = _ans_57_leadingZeros_T_93[23] ? 6'h17 : _ans_57_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_168 = _ans_57_leadingZeros_T_93[22] ? 6'h16 : _ans_57_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_169 = _ans_57_leadingZeros_T_93[21] ? 6'h15 : _ans_57_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_170 = _ans_57_leadingZeros_T_93[20] ? 6'h14 : _ans_57_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_171 = _ans_57_leadingZeros_T_93[19] ? 6'h13 : _ans_57_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_172 = _ans_57_leadingZeros_T_93[18] ? 6'h12 : _ans_57_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_173 = _ans_57_leadingZeros_T_93[17] ? 6'h11 : _ans_57_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_174 = _ans_57_leadingZeros_T_93[16] ? 6'h10 : _ans_57_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_175 = _ans_57_leadingZeros_T_93[15] ? 6'hf : _ans_57_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_176 = _ans_57_leadingZeros_T_93[14] ? 6'he : _ans_57_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_177 = _ans_57_leadingZeros_T_93[13] ? 6'hd : _ans_57_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_178 = _ans_57_leadingZeros_T_93[12] ? 6'hc : _ans_57_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_179 = _ans_57_leadingZeros_T_93[11] ? 6'hb : _ans_57_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_180 = _ans_57_leadingZeros_T_93[10] ? 6'ha : _ans_57_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_181 = _ans_57_leadingZeros_T_93[9] ? 6'h9 : _ans_57_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_182 = _ans_57_leadingZeros_T_93[8] ? 6'h8 : _ans_57_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_183 = _ans_57_leadingZeros_T_93[7] ? 6'h7 : _ans_57_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_184 = _ans_57_leadingZeros_T_93[6] ? 6'h6 : _ans_57_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_185 = _ans_57_leadingZeros_T_93[5] ? 6'h5 : _ans_57_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_186 = _ans_57_leadingZeros_T_93[4] ? 6'h4 : _ans_57_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_187 = _ans_57_leadingZeros_T_93[3] ? 6'h3 : _ans_57_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_188 = _ans_57_leadingZeros_T_93[2] ? 6'h2 : _ans_57_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_leadingZeros_T_189 = _ans_57_leadingZeros_T_93[1] ? 6'h1 : _ans_57_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_57_leadingZeros = _ans_57_leadingZeros_T_93[0] ? 6'h0 : _ans_57_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_57_expRaw_T_1 = 6'h1f - ans_57_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_57_expRaw = ans_57_isZero ? 6'h0 : _ans_57_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_57_shiftAmt_T_2 = ans_57_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_57_shiftAmt = ans_57_expRaw > 6'h3 ? _ans_57_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_57_mantissaRaw_T = ans_57_absClipped >> ans_57_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_57_mantissaRaw = _ans_57_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_57_mantissa = ans_57_expRaw >= 6'h3 ? ans_57_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_57_expAdjusted = ans_57_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_57_exp_T_4 = ans_57_expAdjusted > 7'hf ? 4'hf : ans_57_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_57_exp = ans_57_isZero ? 4'h0 : _ans_57_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_57_fp8 = {ans_57_clippedX[31],ans_57_exp,ans_57_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_58 = {24'h0,linear_bias_58}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_58 = tempSum_58 + biasExtended_58; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_58_sign = sum32_58[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_58_absX_T = ~sum32_58; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_58_absX_T_2 = _ans_58_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_58_absX = ans_58_sign ? _ans_58_absX_T_2 : sum32_58; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_58_shiftedX_T_1 = _GEN_10432 - ans_58_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_58_shiftedX_T_3 = ans_58_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_58_shiftedX = ans_58_sign ? _ans_58_shiftedX_T_1 : _ans_58_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_58_scaledX_T_1 = ans_58_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_58_scaledX = _ans_58_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_58_clippedX_T_2 = ans_58_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_58_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_58_clippedX = ans_58_scaledX > 49'h1c0 ? 49'h1c0 : _ans_58_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_58_absClipped_T_1 = ~ans_58_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_58_absClipped_T_3 = _ans_58_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_58_absClipped = ans_58_clippedX[31] ? _ans_58_absClipped_T_3 : ans_58_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_58_isZero = ans_58_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11072 = {{16'd0}, ans_58_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_4 = _GEN_11072 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_6 = {ans_58_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_8 = _ans_58_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_9 = _ans_58_leadingZeros_T_4 | _ans_58_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11073 = {{8'd0}, _ans_58_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_14 = _GEN_11073 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_16 = {_ans_58_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_18 = _ans_58_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_19 = _ans_58_leadingZeros_T_14 | _ans_58_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11074 = {{4'd0}, _ans_58_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_24 = _GEN_11074 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_26 = {_ans_58_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_28 = _ans_58_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_29 = _ans_58_leadingZeros_T_24 | _ans_58_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11075 = {{2'd0}, _ans_58_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_34 = _GEN_11075 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_36 = {_ans_58_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_38 = _ans_58_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_39 = _ans_58_leadingZeros_T_34 | _ans_58_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11076 = {{1'd0}, _ans_58_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_44 = _GEN_11076 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_46 = {_ans_58_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_48 = _ans_58_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_58_leadingZeros_T_49 = _ans_58_leadingZeros_T_44 | _ans_58_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11077 = {{8'd0}, ans_58_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_55 = _GEN_11077 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_57 = {ans_58_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_59 = _ans_58_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_60 = _ans_58_leadingZeros_T_55 | _ans_58_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11078 = {{4'd0}, _ans_58_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_65 = _GEN_11078 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_67 = {_ans_58_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_69 = _ans_58_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_70 = _ans_58_leadingZeros_T_65 | _ans_58_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11079 = {{2'd0}, _ans_58_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_75 = _GEN_11079 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_77 = {_ans_58_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_79 = _ans_58_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_80 = _ans_58_leadingZeros_T_75 | _ans_58_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11080 = {{1'd0}, _ans_58_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_85 = _GEN_11080 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_87 = {_ans_58_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_89 = _ans_58_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_58_leadingZeros_T_90 = _ans_58_leadingZeros_T_85 | _ans_58_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_58_leadingZeros_T_93 = {_ans_58_leadingZeros_T_49,_ans_58_leadingZeros_T_90,ans_58_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_58_leadingZeros_T_143 = _ans_58_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_144 = _ans_58_leadingZeros_T_93[46] ? 6'h2e : _ans_58_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_145 = _ans_58_leadingZeros_T_93[45] ? 6'h2d : _ans_58_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_146 = _ans_58_leadingZeros_T_93[44] ? 6'h2c : _ans_58_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_147 = _ans_58_leadingZeros_T_93[43] ? 6'h2b : _ans_58_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_148 = _ans_58_leadingZeros_T_93[42] ? 6'h2a : _ans_58_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_149 = _ans_58_leadingZeros_T_93[41] ? 6'h29 : _ans_58_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_150 = _ans_58_leadingZeros_T_93[40] ? 6'h28 : _ans_58_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_151 = _ans_58_leadingZeros_T_93[39] ? 6'h27 : _ans_58_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_152 = _ans_58_leadingZeros_T_93[38] ? 6'h26 : _ans_58_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_153 = _ans_58_leadingZeros_T_93[37] ? 6'h25 : _ans_58_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_154 = _ans_58_leadingZeros_T_93[36] ? 6'h24 : _ans_58_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_155 = _ans_58_leadingZeros_T_93[35] ? 6'h23 : _ans_58_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_156 = _ans_58_leadingZeros_T_93[34] ? 6'h22 : _ans_58_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_157 = _ans_58_leadingZeros_T_93[33] ? 6'h21 : _ans_58_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_158 = _ans_58_leadingZeros_T_93[32] ? 6'h20 : _ans_58_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_159 = _ans_58_leadingZeros_T_93[31] ? 6'h1f : _ans_58_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_160 = _ans_58_leadingZeros_T_93[30] ? 6'h1e : _ans_58_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_161 = _ans_58_leadingZeros_T_93[29] ? 6'h1d : _ans_58_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_162 = _ans_58_leadingZeros_T_93[28] ? 6'h1c : _ans_58_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_163 = _ans_58_leadingZeros_T_93[27] ? 6'h1b : _ans_58_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_164 = _ans_58_leadingZeros_T_93[26] ? 6'h1a : _ans_58_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_165 = _ans_58_leadingZeros_T_93[25] ? 6'h19 : _ans_58_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_166 = _ans_58_leadingZeros_T_93[24] ? 6'h18 : _ans_58_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_167 = _ans_58_leadingZeros_T_93[23] ? 6'h17 : _ans_58_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_168 = _ans_58_leadingZeros_T_93[22] ? 6'h16 : _ans_58_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_169 = _ans_58_leadingZeros_T_93[21] ? 6'h15 : _ans_58_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_170 = _ans_58_leadingZeros_T_93[20] ? 6'h14 : _ans_58_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_171 = _ans_58_leadingZeros_T_93[19] ? 6'h13 : _ans_58_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_172 = _ans_58_leadingZeros_T_93[18] ? 6'h12 : _ans_58_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_173 = _ans_58_leadingZeros_T_93[17] ? 6'h11 : _ans_58_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_174 = _ans_58_leadingZeros_T_93[16] ? 6'h10 : _ans_58_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_175 = _ans_58_leadingZeros_T_93[15] ? 6'hf : _ans_58_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_176 = _ans_58_leadingZeros_T_93[14] ? 6'he : _ans_58_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_177 = _ans_58_leadingZeros_T_93[13] ? 6'hd : _ans_58_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_178 = _ans_58_leadingZeros_T_93[12] ? 6'hc : _ans_58_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_179 = _ans_58_leadingZeros_T_93[11] ? 6'hb : _ans_58_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_180 = _ans_58_leadingZeros_T_93[10] ? 6'ha : _ans_58_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_181 = _ans_58_leadingZeros_T_93[9] ? 6'h9 : _ans_58_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_182 = _ans_58_leadingZeros_T_93[8] ? 6'h8 : _ans_58_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_183 = _ans_58_leadingZeros_T_93[7] ? 6'h7 : _ans_58_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_184 = _ans_58_leadingZeros_T_93[6] ? 6'h6 : _ans_58_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_185 = _ans_58_leadingZeros_T_93[5] ? 6'h5 : _ans_58_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_186 = _ans_58_leadingZeros_T_93[4] ? 6'h4 : _ans_58_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_187 = _ans_58_leadingZeros_T_93[3] ? 6'h3 : _ans_58_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_188 = _ans_58_leadingZeros_T_93[2] ? 6'h2 : _ans_58_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_leadingZeros_T_189 = _ans_58_leadingZeros_T_93[1] ? 6'h1 : _ans_58_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_58_leadingZeros = _ans_58_leadingZeros_T_93[0] ? 6'h0 : _ans_58_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_58_expRaw_T_1 = 6'h1f - ans_58_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_58_expRaw = ans_58_isZero ? 6'h0 : _ans_58_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_58_shiftAmt_T_2 = ans_58_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_58_shiftAmt = ans_58_expRaw > 6'h3 ? _ans_58_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_58_mantissaRaw_T = ans_58_absClipped >> ans_58_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_58_mantissaRaw = _ans_58_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_58_mantissa = ans_58_expRaw >= 6'h3 ? ans_58_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_58_expAdjusted = ans_58_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_58_exp_T_4 = ans_58_expAdjusted > 7'hf ? 4'hf : ans_58_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_58_exp = ans_58_isZero ? 4'h0 : _ans_58_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_58_fp8 = {ans_58_clippedX[31],ans_58_exp,ans_58_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_59 = {24'h0,linear_bias_59}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_59 = tempSum_59 + biasExtended_59; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_59_sign = sum32_59[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_59_absX_T = ~sum32_59; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_59_absX_T_2 = _ans_59_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_59_absX = ans_59_sign ? _ans_59_absX_T_2 : sum32_59; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_59_shiftedX_T_1 = _GEN_10432 - ans_59_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_59_shiftedX_T_3 = ans_59_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_59_shiftedX = ans_59_sign ? _ans_59_shiftedX_T_1 : _ans_59_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_59_scaledX_T_1 = ans_59_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_59_scaledX = _ans_59_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_59_clippedX_T_2 = ans_59_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_59_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_59_clippedX = ans_59_scaledX > 49'h1c0 ? 49'h1c0 : _ans_59_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_59_absClipped_T_1 = ~ans_59_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_59_absClipped_T_3 = _ans_59_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_59_absClipped = ans_59_clippedX[31] ? _ans_59_absClipped_T_3 : ans_59_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_59_isZero = ans_59_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11083 = {{16'd0}, ans_59_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_4 = _GEN_11083 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_6 = {ans_59_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_8 = _ans_59_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_9 = _ans_59_leadingZeros_T_4 | _ans_59_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11084 = {{8'd0}, _ans_59_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_14 = _GEN_11084 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_16 = {_ans_59_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_18 = _ans_59_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_19 = _ans_59_leadingZeros_T_14 | _ans_59_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11085 = {{4'd0}, _ans_59_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_24 = _GEN_11085 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_26 = {_ans_59_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_28 = _ans_59_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_29 = _ans_59_leadingZeros_T_24 | _ans_59_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11086 = {{2'd0}, _ans_59_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_34 = _GEN_11086 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_36 = {_ans_59_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_38 = _ans_59_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_39 = _ans_59_leadingZeros_T_34 | _ans_59_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11087 = {{1'd0}, _ans_59_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_44 = _GEN_11087 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_46 = {_ans_59_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_48 = _ans_59_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_59_leadingZeros_T_49 = _ans_59_leadingZeros_T_44 | _ans_59_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11088 = {{8'd0}, ans_59_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_55 = _GEN_11088 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_57 = {ans_59_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_59 = _ans_59_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_60 = _ans_59_leadingZeros_T_55 | _ans_59_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11089 = {{4'd0}, _ans_59_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_65 = _GEN_11089 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_67 = {_ans_59_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_69 = _ans_59_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_70 = _ans_59_leadingZeros_T_65 | _ans_59_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11090 = {{2'd0}, _ans_59_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_75 = _GEN_11090 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_77 = {_ans_59_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_79 = _ans_59_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_80 = _ans_59_leadingZeros_T_75 | _ans_59_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11091 = {{1'd0}, _ans_59_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_85 = _GEN_11091 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_87 = {_ans_59_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_89 = _ans_59_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_59_leadingZeros_T_90 = _ans_59_leadingZeros_T_85 | _ans_59_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_59_leadingZeros_T_93 = {_ans_59_leadingZeros_T_49,_ans_59_leadingZeros_T_90,ans_59_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_59_leadingZeros_T_143 = _ans_59_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_144 = _ans_59_leadingZeros_T_93[46] ? 6'h2e : _ans_59_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_145 = _ans_59_leadingZeros_T_93[45] ? 6'h2d : _ans_59_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_146 = _ans_59_leadingZeros_T_93[44] ? 6'h2c : _ans_59_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_147 = _ans_59_leadingZeros_T_93[43] ? 6'h2b : _ans_59_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_148 = _ans_59_leadingZeros_T_93[42] ? 6'h2a : _ans_59_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_149 = _ans_59_leadingZeros_T_93[41] ? 6'h29 : _ans_59_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_150 = _ans_59_leadingZeros_T_93[40] ? 6'h28 : _ans_59_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_151 = _ans_59_leadingZeros_T_93[39] ? 6'h27 : _ans_59_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_152 = _ans_59_leadingZeros_T_93[38] ? 6'h26 : _ans_59_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_153 = _ans_59_leadingZeros_T_93[37] ? 6'h25 : _ans_59_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_154 = _ans_59_leadingZeros_T_93[36] ? 6'h24 : _ans_59_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_155 = _ans_59_leadingZeros_T_93[35] ? 6'h23 : _ans_59_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_156 = _ans_59_leadingZeros_T_93[34] ? 6'h22 : _ans_59_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_157 = _ans_59_leadingZeros_T_93[33] ? 6'h21 : _ans_59_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_158 = _ans_59_leadingZeros_T_93[32] ? 6'h20 : _ans_59_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_159 = _ans_59_leadingZeros_T_93[31] ? 6'h1f : _ans_59_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_160 = _ans_59_leadingZeros_T_93[30] ? 6'h1e : _ans_59_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_161 = _ans_59_leadingZeros_T_93[29] ? 6'h1d : _ans_59_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_162 = _ans_59_leadingZeros_T_93[28] ? 6'h1c : _ans_59_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_163 = _ans_59_leadingZeros_T_93[27] ? 6'h1b : _ans_59_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_164 = _ans_59_leadingZeros_T_93[26] ? 6'h1a : _ans_59_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_165 = _ans_59_leadingZeros_T_93[25] ? 6'h19 : _ans_59_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_166 = _ans_59_leadingZeros_T_93[24] ? 6'h18 : _ans_59_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_167 = _ans_59_leadingZeros_T_93[23] ? 6'h17 : _ans_59_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_168 = _ans_59_leadingZeros_T_93[22] ? 6'h16 : _ans_59_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_169 = _ans_59_leadingZeros_T_93[21] ? 6'h15 : _ans_59_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_170 = _ans_59_leadingZeros_T_93[20] ? 6'h14 : _ans_59_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_171 = _ans_59_leadingZeros_T_93[19] ? 6'h13 : _ans_59_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_172 = _ans_59_leadingZeros_T_93[18] ? 6'h12 : _ans_59_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_173 = _ans_59_leadingZeros_T_93[17] ? 6'h11 : _ans_59_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_174 = _ans_59_leadingZeros_T_93[16] ? 6'h10 : _ans_59_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_175 = _ans_59_leadingZeros_T_93[15] ? 6'hf : _ans_59_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_176 = _ans_59_leadingZeros_T_93[14] ? 6'he : _ans_59_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_177 = _ans_59_leadingZeros_T_93[13] ? 6'hd : _ans_59_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_178 = _ans_59_leadingZeros_T_93[12] ? 6'hc : _ans_59_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_179 = _ans_59_leadingZeros_T_93[11] ? 6'hb : _ans_59_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_180 = _ans_59_leadingZeros_T_93[10] ? 6'ha : _ans_59_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_181 = _ans_59_leadingZeros_T_93[9] ? 6'h9 : _ans_59_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_182 = _ans_59_leadingZeros_T_93[8] ? 6'h8 : _ans_59_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_183 = _ans_59_leadingZeros_T_93[7] ? 6'h7 : _ans_59_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_184 = _ans_59_leadingZeros_T_93[6] ? 6'h6 : _ans_59_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_185 = _ans_59_leadingZeros_T_93[5] ? 6'h5 : _ans_59_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_186 = _ans_59_leadingZeros_T_93[4] ? 6'h4 : _ans_59_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_187 = _ans_59_leadingZeros_T_93[3] ? 6'h3 : _ans_59_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_188 = _ans_59_leadingZeros_T_93[2] ? 6'h2 : _ans_59_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_leadingZeros_T_189 = _ans_59_leadingZeros_T_93[1] ? 6'h1 : _ans_59_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_59_leadingZeros = _ans_59_leadingZeros_T_93[0] ? 6'h0 : _ans_59_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_59_expRaw_T_1 = 6'h1f - ans_59_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_59_expRaw = ans_59_isZero ? 6'h0 : _ans_59_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_59_shiftAmt_T_2 = ans_59_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_59_shiftAmt = ans_59_expRaw > 6'h3 ? _ans_59_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_59_mantissaRaw_T = ans_59_absClipped >> ans_59_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_59_mantissaRaw = _ans_59_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_59_mantissa = ans_59_expRaw >= 6'h3 ? ans_59_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_59_expAdjusted = ans_59_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_59_exp_T_4 = ans_59_expAdjusted > 7'hf ? 4'hf : ans_59_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_59_exp = ans_59_isZero ? 4'h0 : _ans_59_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_59_fp8 = {ans_59_clippedX[31],ans_59_exp,ans_59_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_60 = {24'h0,linear_bias_60}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_60 = tempSum_60 + biasExtended_60; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_60_sign = sum32_60[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_60_absX_T = ~sum32_60; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_60_absX_T_2 = _ans_60_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_60_absX = ans_60_sign ? _ans_60_absX_T_2 : sum32_60; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_60_shiftedX_T_1 = _GEN_10432 - ans_60_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_60_shiftedX_T_3 = ans_60_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_60_shiftedX = ans_60_sign ? _ans_60_shiftedX_T_1 : _ans_60_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_60_scaledX_T_1 = ans_60_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_60_scaledX = _ans_60_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_60_clippedX_T_2 = ans_60_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_60_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_60_clippedX = ans_60_scaledX > 49'h1c0 ? 49'h1c0 : _ans_60_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_60_absClipped_T_1 = ~ans_60_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_60_absClipped_T_3 = _ans_60_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_60_absClipped = ans_60_clippedX[31] ? _ans_60_absClipped_T_3 : ans_60_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_60_isZero = ans_60_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11094 = {{16'd0}, ans_60_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_4 = _GEN_11094 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_6 = {ans_60_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_8 = _ans_60_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_9 = _ans_60_leadingZeros_T_4 | _ans_60_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11095 = {{8'd0}, _ans_60_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_14 = _GEN_11095 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_16 = {_ans_60_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_18 = _ans_60_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_19 = _ans_60_leadingZeros_T_14 | _ans_60_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11096 = {{4'd0}, _ans_60_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_24 = _GEN_11096 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_26 = {_ans_60_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_28 = _ans_60_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_29 = _ans_60_leadingZeros_T_24 | _ans_60_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11097 = {{2'd0}, _ans_60_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_34 = _GEN_11097 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_36 = {_ans_60_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_38 = _ans_60_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_39 = _ans_60_leadingZeros_T_34 | _ans_60_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11098 = {{1'd0}, _ans_60_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_44 = _GEN_11098 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_46 = {_ans_60_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_48 = _ans_60_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_60_leadingZeros_T_49 = _ans_60_leadingZeros_T_44 | _ans_60_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11099 = {{8'd0}, ans_60_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_55 = _GEN_11099 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_57 = {ans_60_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_59 = _ans_60_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_60 = _ans_60_leadingZeros_T_55 | _ans_60_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11100 = {{4'd0}, _ans_60_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_65 = _GEN_11100 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_67 = {_ans_60_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_69 = _ans_60_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_70 = _ans_60_leadingZeros_T_65 | _ans_60_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11101 = {{2'd0}, _ans_60_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_75 = _GEN_11101 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_77 = {_ans_60_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_79 = _ans_60_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_80 = _ans_60_leadingZeros_T_75 | _ans_60_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11102 = {{1'd0}, _ans_60_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_85 = _GEN_11102 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_87 = {_ans_60_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_89 = _ans_60_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_60_leadingZeros_T_90 = _ans_60_leadingZeros_T_85 | _ans_60_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_60_leadingZeros_T_93 = {_ans_60_leadingZeros_T_49,_ans_60_leadingZeros_T_90,ans_60_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_60_leadingZeros_T_143 = _ans_60_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_144 = _ans_60_leadingZeros_T_93[46] ? 6'h2e : _ans_60_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_145 = _ans_60_leadingZeros_T_93[45] ? 6'h2d : _ans_60_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_146 = _ans_60_leadingZeros_T_93[44] ? 6'h2c : _ans_60_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_147 = _ans_60_leadingZeros_T_93[43] ? 6'h2b : _ans_60_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_148 = _ans_60_leadingZeros_T_93[42] ? 6'h2a : _ans_60_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_149 = _ans_60_leadingZeros_T_93[41] ? 6'h29 : _ans_60_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_150 = _ans_60_leadingZeros_T_93[40] ? 6'h28 : _ans_60_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_151 = _ans_60_leadingZeros_T_93[39] ? 6'h27 : _ans_60_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_152 = _ans_60_leadingZeros_T_93[38] ? 6'h26 : _ans_60_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_153 = _ans_60_leadingZeros_T_93[37] ? 6'h25 : _ans_60_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_154 = _ans_60_leadingZeros_T_93[36] ? 6'h24 : _ans_60_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_155 = _ans_60_leadingZeros_T_93[35] ? 6'h23 : _ans_60_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_156 = _ans_60_leadingZeros_T_93[34] ? 6'h22 : _ans_60_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_157 = _ans_60_leadingZeros_T_93[33] ? 6'h21 : _ans_60_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_158 = _ans_60_leadingZeros_T_93[32] ? 6'h20 : _ans_60_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_159 = _ans_60_leadingZeros_T_93[31] ? 6'h1f : _ans_60_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_160 = _ans_60_leadingZeros_T_93[30] ? 6'h1e : _ans_60_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_161 = _ans_60_leadingZeros_T_93[29] ? 6'h1d : _ans_60_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_162 = _ans_60_leadingZeros_T_93[28] ? 6'h1c : _ans_60_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_163 = _ans_60_leadingZeros_T_93[27] ? 6'h1b : _ans_60_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_164 = _ans_60_leadingZeros_T_93[26] ? 6'h1a : _ans_60_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_165 = _ans_60_leadingZeros_T_93[25] ? 6'h19 : _ans_60_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_166 = _ans_60_leadingZeros_T_93[24] ? 6'h18 : _ans_60_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_167 = _ans_60_leadingZeros_T_93[23] ? 6'h17 : _ans_60_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_168 = _ans_60_leadingZeros_T_93[22] ? 6'h16 : _ans_60_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_169 = _ans_60_leadingZeros_T_93[21] ? 6'h15 : _ans_60_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_170 = _ans_60_leadingZeros_T_93[20] ? 6'h14 : _ans_60_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_171 = _ans_60_leadingZeros_T_93[19] ? 6'h13 : _ans_60_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_172 = _ans_60_leadingZeros_T_93[18] ? 6'h12 : _ans_60_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_173 = _ans_60_leadingZeros_T_93[17] ? 6'h11 : _ans_60_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_174 = _ans_60_leadingZeros_T_93[16] ? 6'h10 : _ans_60_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_175 = _ans_60_leadingZeros_T_93[15] ? 6'hf : _ans_60_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_176 = _ans_60_leadingZeros_T_93[14] ? 6'he : _ans_60_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_177 = _ans_60_leadingZeros_T_93[13] ? 6'hd : _ans_60_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_178 = _ans_60_leadingZeros_T_93[12] ? 6'hc : _ans_60_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_179 = _ans_60_leadingZeros_T_93[11] ? 6'hb : _ans_60_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_180 = _ans_60_leadingZeros_T_93[10] ? 6'ha : _ans_60_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_181 = _ans_60_leadingZeros_T_93[9] ? 6'h9 : _ans_60_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_182 = _ans_60_leadingZeros_T_93[8] ? 6'h8 : _ans_60_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_183 = _ans_60_leadingZeros_T_93[7] ? 6'h7 : _ans_60_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_184 = _ans_60_leadingZeros_T_93[6] ? 6'h6 : _ans_60_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_185 = _ans_60_leadingZeros_T_93[5] ? 6'h5 : _ans_60_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_186 = _ans_60_leadingZeros_T_93[4] ? 6'h4 : _ans_60_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_187 = _ans_60_leadingZeros_T_93[3] ? 6'h3 : _ans_60_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_188 = _ans_60_leadingZeros_T_93[2] ? 6'h2 : _ans_60_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_leadingZeros_T_189 = _ans_60_leadingZeros_T_93[1] ? 6'h1 : _ans_60_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_60_leadingZeros = _ans_60_leadingZeros_T_93[0] ? 6'h0 : _ans_60_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_60_expRaw_T_1 = 6'h1f - ans_60_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_60_expRaw = ans_60_isZero ? 6'h0 : _ans_60_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_60_shiftAmt_T_2 = ans_60_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_60_shiftAmt = ans_60_expRaw > 6'h3 ? _ans_60_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_60_mantissaRaw_T = ans_60_absClipped >> ans_60_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_60_mantissaRaw = _ans_60_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_60_mantissa = ans_60_expRaw >= 6'h3 ? ans_60_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_60_expAdjusted = ans_60_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_60_exp_T_4 = ans_60_expAdjusted > 7'hf ? 4'hf : ans_60_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_60_exp = ans_60_isZero ? 4'h0 : _ans_60_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_60_fp8 = {ans_60_clippedX[31],ans_60_exp,ans_60_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_61 = {24'h0,linear_bias_61}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_61 = tempSum_61 + biasExtended_61; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_61_sign = sum32_61[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_61_absX_T = ~sum32_61; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_61_absX_T_2 = _ans_61_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_61_absX = ans_61_sign ? _ans_61_absX_T_2 : sum32_61; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_61_shiftedX_T_1 = _GEN_10432 - ans_61_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_61_shiftedX_T_3 = ans_61_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_61_shiftedX = ans_61_sign ? _ans_61_shiftedX_T_1 : _ans_61_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_61_scaledX_T_1 = ans_61_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_61_scaledX = _ans_61_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_61_clippedX_T_2 = ans_61_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_61_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_61_clippedX = ans_61_scaledX > 49'h1c0 ? 49'h1c0 : _ans_61_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_61_absClipped_T_1 = ~ans_61_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_61_absClipped_T_3 = _ans_61_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_61_absClipped = ans_61_clippedX[31] ? _ans_61_absClipped_T_3 : ans_61_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_61_isZero = ans_61_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11105 = {{16'd0}, ans_61_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_4 = _GEN_11105 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_6 = {ans_61_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_8 = _ans_61_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_9 = _ans_61_leadingZeros_T_4 | _ans_61_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11106 = {{8'd0}, _ans_61_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_14 = _GEN_11106 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_16 = {_ans_61_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_18 = _ans_61_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_19 = _ans_61_leadingZeros_T_14 | _ans_61_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11107 = {{4'd0}, _ans_61_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_24 = _GEN_11107 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_26 = {_ans_61_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_28 = _ans_61_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_29 = _ans_61_leadingZeros_T_24 | _ans_61_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11108 = {{2'd0}, _ans_61_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_34 = _GEN_11108 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_36 = {_ans_61_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_38 = _ans_61_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_39 = _ans_61_leadingZeros_T_34 | _ans_61_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11109 = {{1'd0}, _ans_61_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_44 = _GEN_11109 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_46 = {_ans_61_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_48 = _ans_61_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_61_leadingZeros_T_49 = _ans_61_leadingZeros_T_44 | _ans_61_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11110 = {{8'd0}, ans_61_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_55 = _GEN_11110 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_57 = {ans_61_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_59 = _ans_61_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_60 = _ans_61_leadingZeros_T_55 | _ans_61_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11111 = {{4'd0}, _ans_61_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_65 = _GEN_11111 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_67 = {_ans_61_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_69 = _ans_61_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_70 = _ans_61_leadingZeros_T_65 | _ans_61_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11112 = {{2'd0}, _ans_61_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_75 = _GEN_11112 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_77 = {_ans_61_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_79 = _ans_61_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_80 = _ans_61_leadingZeros_T_75 | _ans_61_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11113 = {{1'd0}, _ans_61_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_85 = _GEN_11113 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_87 = {_ans_61_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_89 = _ans_61_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_61_leadingZeros_T_90 = _ans_61_leadingZeros_T_85 | _ans_61_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_61_leadingZeros_T_93 = {_ans_61_leadingZeros_T_49,_ans_61_leadingZeros_T_90,ans_61_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_61_leadingZeros_T_143 = _ans_61_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_144 = _ans_61_leadingZeros_T_93[46] ? 6'h2e : _ans_61_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_145 = _ans_61_leadingZeros_T_93[45] ? 6'h2d : _ans_61_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_146 = _ans_61_leadingZeros_T_93[44] ? 6'h2c : _ans_61_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_147 = _ans_61_leadingZeros_T_93[43] ? 6'h2b : _ans_61_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_148 = _ans_61_leadingZeros_T_93[42] ? 6'h2a : _ans_61_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_149 = _ans_61_leadingZeros_T_93[41] ? 6'h29 : _ans_61_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_150 = _ans_61_leadingZeros_T_93[40] ? 6'h28 : _ans_61_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_151 = _ans_61_leadingZeros_T_93[39] ? 6'h27 : _ans_61_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_152 = _ans_61_leadingZeros_T_93[38] ? 6'h26 : _ans_61_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_153 = _ans_61_leadingZeros_T_93[37] ? 6'h25 : _ans_61_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_154 = _ans_61_leadingZeros_T_93[36] ? 6'h24 : _ans_61_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_155 = _ans_61_leadingZeros_T_93[35] ? 6'h23 : _ans_61_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_156 = _ans_61_leadingZeros_T_93[34] ? 6'h22 : _ans_61_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_157 = _ans_61_leadingZeros_T_93[33] ? 6'h21 : _ans_61_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_158 = _ans_61_leadingZeros_T_93[32] ? 6'h20 : _ans_61_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_159 = _ans_61_leadingZeros_T_93[31] ? 6'h1f : _ans_61_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_160 = _ans_61_leadingZeros_T_93[30] ? 6'h1e : _ans_61_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_161 = _ans_61_leadingZeros_T_93[29] ? 6'h1d : _ans_61_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_162 = _ans_61_leadingZeros_T_93[28] ? 6'h1c : _ans_61_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_163 = _ans_61_leadingZeros_T_93[27] ? 6'h1b : _ans_61_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_164 = _ans_61_leadingZeros_T_93[26] ? 6'h1a : _ans_61_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_165 = _ans_61_leadingZeros_T_93[25] ? 6'h19 : _ans_61_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_166 = _ans_61_leadingZeros_T_93[24] ? 6'h18 : _ans_61_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_167 = _ans_61_leadingZeros_T_93[23] ? 6'h17 : _ans_61_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_168 = _ans_61_leadingZeros_T_93[22] ? 6'h16 : _ans_61_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_169 = _ans_61_leadingZeros_T_93[21] ? 6'h15 : _ans_61_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_170 = _ans_61_leadingZeros_T_93[20] ? 6'h14 : _ans_61_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_171 = _ans_61_leadingZeros_T_93[19] ? 6'h13 : _ans_61_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_172 = _ans_61_leadingZeros_T_93[18] ? 6'h12 : _ans_61_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_173 = _ans_61_leadingZeros_T_93[17] ? 6'h11 : _ans_61_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_174 = _ans_61_leadingZeros_T_93[16] ? 6'h10 : _ans_61_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_175 = _ans_61_leadingZeros_T_93[15] ? 6'hf : _ans_61_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_176 = _ans_61_leadingZeros_T_93[14] ? 6'he : _ans_61_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_177 = _ans_61_leadingZeros_T_93[13] ? 6'hd : _ans_61_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_178 = _ans_61_leadingZeros_T_93[12] ? 6'hc : _ans_61_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_179 = _ans_61_leadingZeros_T_93[11] ? 6'hb : _ans_61_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_180 = _ans_61_leadingZeros_T_93[10] ? 6'ha : _ans_61_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_181 = _ans_61_leadingZeros_T_93[9] ? 6'h9 : _ans_61_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_182 = _ans_61_leadingZeros_T_93[8] ? 6'h8 : _ans_61_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_183 = _ans_61_leadingZeros_T_93[7] ? 6'h7 : _ans_61_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_184 = _ans_61_leadingZeros_T_93[6] ? 6'h6 : _ans_61_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_185 = _ans_61_leadingZeros_T_93[5] ? 6'h5 : _ans_61_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_186 = _ans_61_leadingZeros_T_93[4] ? 6'h4 : _ans_61_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_187 = _ans_61_leadingZeros_T_93[3] ? 6'h3 : _ans_61_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_188 = _ans_61_leadingZeros_T_93[2] ? 6'h2 : _ans_61_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_leadingZeros_T_189 = _ans_61_leadingZeros_T_93[1] ? 6'h1 : _ans_61_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_61_leadingZeros = _ans_61_leadingZeros_T_93[0] ? 6'h0 : _ans_61_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_61_expRaw_T_1 = 6'h1f - ans_61_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_61_expRaw = ans_61_isZero ? 6'h0 : _ans_61_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_61_shiftAmt_T_2 = ans_61_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_61_shiftAmt = ans_61_expRaw > 6'h3 ? _ans_61_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_61_mantissaRaw_T = ans_61_absClipped >> ans_61_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_61_mantissaRaw = _ans_61_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_61_mantissa = ans_61_expRaw >= 6'h3 ? ans_61_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_61_expAdjusted = ans_61_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_61_exp_T_4 = ans_61_expAdjusted > 7'hf ? 4'hf : ans_61_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_61_exp = ans_61_isZero ? 4'h0 : _ans_61_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_61_fp8 = {ans_61_clippedX[31],ans_61_exp,ans_61_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_62 = {24'h0,linear_bias_62}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_62 = tempSum_62 + biasExtended_62; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_62_sign = sum32_62[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_62_absX_T = ~sum32_62; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_62_absX_T_2 = _ans_62_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_62_absX = ans_62_sign ? _ans_62_absX_T_2 : sum32_62; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_62_shiftedX_T_1 = _GEN_10432 - ans_62_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_62_shiftedX_T_3 = ans_62_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_62_shiftedX = ans_62_sign ? _ans_62_shiftedX_T_1 : _ans_62_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_62_scaledX_T_1 = ans_62_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_62_scaledX = _ans_62_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_62_clippedX_T_2 = ans_62_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_62_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_62_clippedX = ans_62_scaledX > 49'h1c0 ? 49'h1c0 : _ans_62_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_62_absClipped_T_1 = ~ans_62_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_62_absClipped_T_3 = _ans_62_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_62_absClipped = ans_62_clippedX[31] ? _ans_62_absClipped_T_3 : ans_62_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_62_isZero = ans_62_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11116 = {{16'd0}, ans_62_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_4 = _GEN_11116 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_6 = {ans_62_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_8 = _ans_62_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_9 = _ans_62_leadingZeros_T_4 | _ans_62_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11117 = {{8'd0}, _ans_62_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_14 = _GEN_11117 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_16 = {_ans_62_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_18 = _ans_62_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_19 = _ans_62_leadingZeros_T_14 | _ans_62_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11118 = {{4'd0}, _ans_62_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_24 = _GEN_11118 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_26 = {_ans_62_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_28 = _ans_62_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_29 = _ans_62_leadingZeros_T_24 | _ans_62_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11119 = {{2'd0}, _ans_62_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_34 = _GEN_11119 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_36 = {_ans_62_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_38 = _ans_62_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_39 = _ans_62_leadingZeros_T_34 | _ans_62_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11120 = {{1'd0}, _ans_62_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_44 = _GEN_11120 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_46 = {_ans_62_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_48 = _ans_62_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_62_leadingZeros_T_49 = _ans_62_leadingZeros_T_44 | _ans_62_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11121 = {{8'd0}, ans_62_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_55 = _GEN_11121 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_57 = {ans_62_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_59 = _ans_62_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_60 = _ans_62_leadingZeros_T_55 | _ans_62_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11122 = {{4'd0}, _ans_62_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_65 = _GEN_11122 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_67 = {_ans_62_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_69 = _ans_62_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_70 = _ans_62_leadingZeros_T_65 | _ans_62_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11123 = {{2'd0}, _ans_62_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_75 = _GEN_11123 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_77 = {_ans_62_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_79 = _ans_62_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_80 = _ans_62_leadingZeros_T_75 | _ans_62_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11124 = {{1'd0}, _ans_62_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_85 = _GEN_11124 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_87 = {_ans_62_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_89 = _ans_62_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_62_leadingZeros_T_90 = _ans_62_leadingZeros_T_85 | _ans_62_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_62_leadingZeros_T_93 = {_ans_62_leadingZeros_T_49,_ans_62_leadingZeros_T_90,ans_62_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_62_leadingZeros_T_143 = _ans_62_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_144 = _ans_62_leadingZeros_T_93[46] ? 6'h2e : _ans_62_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_145 = _ans_62_leadingZeros_T_93[45] ? 6'h2d : _ans_62_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_146 = _ans_62_leadingZeros_T_93[44] ? 6'h2c : _ans_62_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_147 = _ans_62_leadingZeros_T_93[43] ? 6'h2b : _ans_62_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_148 = _ans_62_leadingZeros_T_93[42] ? 6'h2a : _ans_62_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_149 = _ans_62_leadingZeros_T_93[41] ? 6'h29 : _ans_62_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_150 = _ans_62_leadingZeros_T_93[40] ? 6'h28 : _ans_62_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_151 = _ans_62_leadingZeros_T_93[39] ? 6'h27 : _ans_62_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_152 = _ans_62_leadingZeros_T_93[38] ? 6'h26 : _ans_62_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_153 = _ans_62_leadingZeros_T_93[37] ? 6'h25 : _ans_62_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_154 = _ans_62_leadingZeros_T_93[36] ? 6'h24 : _ans_62_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_155 = _ans_62_leadingZeros_T_93[35] ? 6'h23 : _ans_62_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_156 = _ans_62_leadingZeros_T_93[34] ? 6'h22 : _ans_62_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_157 = _ans_62_leadingZeros_T_93[33] ? 6'h21 : _ans_62_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_158 = _ans_62_leadingZeros_T_93[32] ? 6'h20 : _ans_62_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_159 = _ans_62_leadingZeros_T_93[31] ? 6'h1f : _ans_62_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_160 = _ans_62_leadingZeros_T_93[30] ? 6'h1e : _ans_62_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_161 = _ans_62_leadingZeros_T_93[29] ? 6'h1d : _ans_62_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_162 = _ans_62_leadingZeros_T_93[28] ? 6'h1c : _ans_62_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_163 = _ans_62_leadingZeros_T_93[27] ? 6'h1b : _ans_62_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_164 = _ans_62_leadingZeros_T_93[26] ? 6'h1a : _ans_62_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_165 = _ans_62_leadingZeros_T_93[25] ? 6'h19 : _ans_62_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_166 = _ans_62_leadingZeros_T_93[24] ? 6'h18 : _ans_62_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_167 = _ans_62_leadingZeros_T_93[23] ? 6'h17 : _ans_62_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_168 = _ans_62_leadingZeros_T_93[22] ? 6'h16 : _ans_62_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_169 = _ans_62_leadingZeros_T_93[21] ? 6'h15 : _ans_62_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_170 = _ans_62_leadingZeros_T_93[20] ? 6'h14 : _ans_62_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_171 = _ans_62_leadingZeros_T_93[19] ? 6'h13 : _ans_62_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_172 = _ans_62_leadingZeros_T_93[18] ? 6'h12 : _ans_62_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_173 = _ans_62_leadingZeros_T_93[17] ? 6'h11 : _ans_62_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_174 = _ans_62_leadingZeros_T_93[16] ? 6'h10 : _ans_62_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_175 = _ans_62_leadingZeros_T_93[15] ? 6'hf : _ans_62_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_176 = _ans_62_leadingZeros_T_93[14] ? 6'he : _ans_62_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_177 = _ans_62_leadingZeros_T_93[13] ? 6'hd : _ans_62_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_178 = _ans_62_leadingZeros_T_93[12] ? 6'hc : _ans_62_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_179 = _ans_62_leadingZeros_T_93[11] ? 6'hb : _ans_62_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_180 = _ans_62_leadingZeros_T_93[10] ? 6'ha : _ans_62_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_181 = _ans_62_leadingZeros_T_93[9] ? 6'h9 : _ans_62_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_182 = _ans_62_leadingZeros_T_93[8] ? 6'h8 : _ans_62_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_183 = _ans_62_leadingZeros_T_93[7] ? 6'h7 : _ans_62_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_184 = _ans_62_leadingZeros_T_93[6] ? 6'h6 : _ans_62_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_185 = _ans_62_leadingZeros_T_93[5] ? 6'h5 : _ans_62_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_186 = _ans_62_leadingZeros_T_93[4] ? 6'h4 : _ans_62_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_187 = _ans_62_leadingZeros_T_93[3] ? 6'h3 : _ans_62_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_188 = _ans_62_leadingZeros_T_93[2] ? 6'h2 : _ans_62_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_leadingZeros_T_189 = _ans_62_leadingZeros_T_93[1] ? 6'h1 : _ans_62_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_62_leadingZeros = _ans_62_leadingZeros_T_93[0] ? 6'h0 : _ans_62_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_62_expRaw_T_1 = 6'h1f - ans_62_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_62_expRaw = ans_62_isZero ? 6'h0 : _ans_62_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_62_shiftAmt_T_2 = ans_62_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_62_shiftAmt = ans_62_expRaw > 6'h3 ? _ans_62_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_62_mantissaRaw_T = ans_62_absClipped >> ans_62_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_62_mantissaRaw = _ans_62_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_62_mantissa = ans_62_expRaw >= 6'h3 ? ans_62_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_62_expAdjusted = ans_62_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_62_exp_T_4 = ans_62_expAdjusted > 7'hf ? 4'hf : ans_62_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_62_exp = ans_62_isZero ? 4'h0 : _ans_62_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_62_fp8 = {ans_62_clippedX[31],ans_62_exp,ans_62_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [31:0] biasExtended_63 = {24'h0,linear_bias_63}; // @[src/main/scala/Multiple/LinearCompute.scala 100:31]
  wire [31:0] sum32_63 = tempSum_63 + biasExtended_63; // @[src/main/scala/Multiple/LinearCompute.scala 101:32]
  wire  ans_63_sign = sum32_63[31]; // @[src/main/scala/Multiple/LinearCompute.scala 37:21]
  wire [31:0] _ans_63_absX_T = ~sum32_63; // @[src/main/scala/Multiple/LinearCompute.scala 38:31]
  wire [31:0] _ans_63_absX_T_2 = _ans_63_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 38:34]
  wire [31:0] ans_63_absX = ans_63_sign ? _ans_63_absX_T_2 : sum32_63; // @[src/main/scala/Multiple/LinearCompute.scala 38:23]
  wire [31:0] _ans_63_shiftedX_T_1 = _GEN_10432 - ans_63_absX; // @[src/main/scala/Multiple/LinearCompute.scala 41:44]
  wire [31:0] _ans_63_shiftedX_T_3 = ans_63_absX - _GEN_10432; // @[src/main/scala/Multiple/LinearCompute.scala 41:57]
  wire [31:0] ans_63_shiftedX = ans_63_sign ? _ans_63_shiftedX_T_1 : _ans_63_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 41:27]
  wire [48:0] _ans_63_scaledX_T_1 = ans_63_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 42:33]
  wire [48:0] ans_63_scaledX = _ans_63_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 42:48]
  wire [48:0] _ans_63_clippedX_T_2 = ans_63_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_63_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 49:59]
  wire [48:0] ans_63_clippedX = ans_63_scaledX > 49'h1c0 ? 49'h1c0 : _ans_63_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 49:27]
  wire [48:0] _ans_63_absClipped_T_1 = ~ans_63_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:45]
  wire [48:0] _ans_63_absClipped_T_3 = _ans_63_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 52:55]
  wire [48:0] ans_63_absClipped = ans_63_clippedX[31] ? _ans_63_absClipped_T_3 : ans_63_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 52:29]
  wire  ans_63_isZero = ans_63_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 53:33]
  wire [31:0] _GEN_11127 = {{16'd0}, ans_63_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_4 = _GEN_11127 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_6 = {ans_63_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_8 = _ans_63_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_9 = _ans_63_leadingZeros_T_4 | _ans_63_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11128 = {{8'd0}, _ans_63_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_14 = _GEN_11128 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_16 = {_ans_63_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_18 = _ans_63_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_19 = _ans_63_leadingZeros_T_14 | _ans_63_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11129 = {{4'd0}, _ans_63_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_24 = _GEN_11129 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_26 = {_ans_63_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_28 = _ans_63_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_29 = _ans_63_leadingZeros_T_24 | _ans_63_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11130 = {{2'd0}, _ans_63_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_34 = _GEN_11130 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_36 = {_ans_63_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_38 = _ans_63_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_39 = _ans_63_leadingZeros_T_34 | _ans_63_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _GEN_11131 = {{1'd0}, _ans_63_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_44 = _GEN_11131 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_46 = {_ans_63_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_48 = _ans_63_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [31:0] _ans_63_leadingZeros_T_49 = _ans_63_leadingZeros_T_44 | _ans_63_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11132 = {{8'd0}, ans_63_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_55 = _GEN_11132 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_57 = {ans_63_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_59 = _ans_63_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_60 = _ans_63_leadingZeros_T_55 | _ans_63_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11133 = {{4'd0}, _ans_63_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_65 = _GEN_11133 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_67 = {_ans_63_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_69 = _ans_63_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_70 = _ans_63_leadingZeros_T_65 | _ans_63_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11134 = {{2'd0}, _ans_63_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_75 = _GEN_11134 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_77 = {_ans_63_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_79 = _ans_63_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_80 = _ans_63_leadingZeros_T_75 | _ans_63_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _GEN_11135 = {{1'd0}, _ans_63_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_85 = _GEN_11135 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_87 = {_ans_63_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_89 = _ans_63_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [15:0] _ans_63_leadingZeros_T_90 = _ans_63_leadingZeros_T_85 | _ans_63_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [48:0] _ans_63_leadingZeros_T_93 = {_ans_63_leadingZeros_T_49,_ans_63_leadingZeros_T_90,ans_63_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 54:51]
  wire [5:0] _ans_63_leadingZeros_T_143 = _ans_63_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_144 = _ans_63_leadingZeros_T_93[46] ? 6'h2e : _ans_63_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_145 = _ans_63_leadingZeros_T_93[45] ? 6'h2d : _ans_63_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_146 = _ans_63_leadingZeros_T_93[44] ? 6'h2c : _ans_63_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_147 = _ans_63_leadingZeros_T_93[43] ? 6'h2b : _ans_63_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_148 = _ans_63_leadingZeros_T_93[42] ? 6'h2a : _ans_63_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_149 = _ans_63_leadingZeros_T_93[41] ? 6'h29 : _ans_63_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_150 = _ans_63_leadingZeros_T_93[40] ? 6'h28 : _ans_63_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_151 = _ans_63_leadingZeros_T_93[39] ? 6'h27 : _ans_63_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_152 = _ans_63_leadingZeros_T_93[38] ? 6'h26 : _ans_63_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_153 = _ans_63_leadingZeros_T_93[37] ? 6'h25 : _ans_63_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_154 = _ans_63_leadingZeros_T_93[36] ? 6'h24 : _ans_63_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_155 = _ans_63_leadingZeros_T_93[35] ? 6'h23 : _ans_63_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_156 = _ans_63_leadingZeros_T_93[34] ? 6'h22 : _ans_63_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_157 = _ans_63_leadingZeros_T_93[33] ? 6'h21 : _ans_63_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_158 = _ans_63_leadingZeros_T_93[32] ? 6'h20 : _ans_63_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_159 = _ans_63_leadingZeros_T_93[31] ? 6'h1f : _ans_63_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_160 = _ans_63_leadingZeros_T_93[30] ? 6'h1e : _ans_63_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_161 = _ans_63_leadingZeros_T_93[29] ? 6'h1d : _ans_63_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_162 = _ans_63_leadingZeros_T_93[28] ? 6'h1c : _ans_63_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_163 = _ans_63_leadingZeros_T_93[27] ? 6'h1b : _ans_63_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_164 = _ans_63_leadingZeros_T_93[26] ? 6'h1a : _ans_63_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_165 = _ans_63_leadingZeros_T_93[25] ? 6'h19 : _ans_63_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_166 = _ans_63_leadingZeros_T_93[24] ? 6'h18 : _ans_63_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_167 = _ans_63_leadingZeros_T_93[23] ? 6'h17 : _ans_63_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_168 = _ans_63_leadingZeros_T_93[22] ? 6'h16 : _ans_63_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_169 = _ans_63_leadingZeros_T_93[21] ? 6'h15 : _ans_63_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_170 = _ans_63_leadingZeros_T_93[20] ? 6'h14 : _ans_63_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_171 = _ans_63_leadingZeros_T_93[19] ? 6'h13 : _ans_63_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_172 = _ans_63_leadingZeros_T_93[18] ? 6'h12 : _ans_63_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_173 = _ans_63_leadingZeros_T_93[17] ? 6'h11 : _ans_63_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_174 = _ans_63_leadingZeros_T_93[16] ? 6'h10 : _ans_63_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_175 = _ans_63_leadingZeros_T_93[15] ? 6'hf : _ans_63_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_176 = _ans_63_leadingZeros_T_93[14] ? 6'he : _ans_63_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_177 = _ans_63_leadingZeros_T_93[13] ? 6'hd : _ans_63_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_178 = _ans_63_leadingZeros_T_93[12] ? 6'hc : _ans_63_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_179 = _ans_63_leadingZeros_T_93[11] ? 6'hb : _ans_63_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_180 = _ans_63_leadingZeros_T_93[10] ? 6'ha : _ans_63_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_181 = _ans_63_leadingZeros_T_93[9] ? 6'h9 : _ans_63_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_182 = _ans_63_leadingZeros_T_93[8] ? 6'h8 : _ans_63_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_183 = _ans_63_leadingZeros_T_93[7] ? 6'h7 : _ans_63_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_184 = _ans_63_leadingZeros_T_93[6] ? 6'h6 : _ans_63_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_185 = _ans_63_leadingZeros_T_93[5] ? 6'h5 : _ans_63_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_186 = _ans_63_leadingZeros_T_93[4] ? 6'h4 : _ans_63_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_187 = _ans_63_leadingZeros_T_93[3] ? 6'h3 : _ans_63_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_188 = _ans_63_leadingZeros_T_93[2] ? 6'h2 : _ans_63_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_leadingZeros_T_189 = _ans_63_leadingZeros_T_93[1] ? 6'h1 : _ans_63_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_63_leadingZeros = _ans_63_leadingZeros_T_93[0] ? 6'h0 : _ans_63_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_63_expRaw_T_1 = 6'h1f - ans_63_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 55:44]
  wire [5:0] ans_63_expRaw = ans_63_isZero ? 6'h0 : _ans_63_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 55:25]
  wire [5:0] _ans_63_shiftAmt_T_2 = ans_63_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 61:49]
  wire [5:0] ans_63_shiftAmt = ans_63_expRaw > 6'h3 ? _ans_63_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 61:27]
  wire [48:0] _ans_63_mantissaRaw_T = ans_63_absClipped >> ans_63_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 62:39]
  wire [6:0] ans_63_mantissaRaw = _ans_63_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 62:51]
  wire [2:0] ans_63_mantissa = ans_63_expRaw >= 6'h3 ? ans_63_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 63:27]
  wire [6:0] ans_63_expAdjusted = ans_63_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 65:34]
  wire [3:0] _ans_63_exp_T_4 = ans_63_expAdjusted > 7'hf ? 4'hf : ans_63_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 66:39]
  wire [3:0] ans_63_exp = ans_63_isZero ? 4'h0 : _ans_63_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 66:22]
  wire [7:0] ans_63_fp8 = {ans_63_clippedX[31],ans_63_exp,ans_63_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 68:22]
  wire [7:0] io_featuresOut_0_scaledX = {{2'd0}, ans_0[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_0_sum = io_featuresOut_0_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_0_minVal = io_featuresOut_0_sum < 8'h40 ? io_featuresOut_0_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_1_scaledX = {{2'd0}, ans_1[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_1_sum = io_featuresOut_1_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_1_minVal = io_featuresOut_1_sum < 8'h40 ? io_featuresOut_1_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_2_scaledX = {{2'd0}, ans_2[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_2_sum = io_featuresOut_2_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_2_minVal = io_featuresOut_2_sum < 8'h40 ? io_featuresOut_2_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_3_scaledX = {{2'd0}, ans_3[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_3_sum = io_featuresOut_3_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_3_minVal = io_featuresOut_3_sum < 8'h40 ? io_featuresOut_3_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_4_scaledX = {{2'd0}, ans_4[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_4_sum = io_featuresOut_4_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_4_minVal = io_featuresOut_4_sum < 8'h40 ? io_featuresOut_4_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_5_scaledX = {{2'd0}, ans_5[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_5_sum = io_featuresOut_5_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_5_minVal = io_featuresOut_5_sum < 8'h40 ? io_featuresOut_5_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_6_scaledX = {{2'd0}, ans_6[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_6_sum = io_featuresOut_6_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_6_minVal = io_featuresOut_6_sum < 8'h40 ? io_featuresOut_6_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_7_scaledX = {{2'd0}, ans_7[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_7_sum = io_featuresOut_7_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_7_minVal = io_featuresOut_7_sum < 8'h40 ? io_featuresOut_7_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_8_scaledX = {{2'd0}, ans_8[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_8_sum = io_featuresOut_8_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_8_minVal = io_featuresOut_8_sum < 8'h40 ? io_featuresOut_8_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_9_scaledX = {{2'd0}, ans_9[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_9_sum = io_featuresOut_9_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_9_minVal = io_featuresOut_9_sum < 8'h40 ? io_featuresOut_9_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_10_scaledX = {{2'd0}, ans_10[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_10_sum = io_featuresOut_10_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_10_minVal = io_featuresOut_10_sum < 8'h40 ? io_featuresOut_10_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_11_scaledX = {{2'd0}, ans_11[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_11_sum = io_featuresOut_11_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_11_minVal = io_featuresOut_11_sum < 8'h40 ? io_featuresOut_11_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_12_scaledX = {{2'd0}, ans_12[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_12_sum = io_featuresOut_12_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_12_minVal = io_featuresOut_12_sum < 8'h40 ? io_featuresOut_12_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_13_scaledX = {{2'd0}, ans_13[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_13_sum = io_featuresOut_13_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_13_minVal = io_featuresOut_13_sum < 8'h40 ? io_featuresOut_13_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_14_scaledX = {{2'd0}, ans_14[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_14_sum = io_featuresOut_14_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_14_minVal = io_featuresOut_14_sum < 8'h40 ? io_featuresOut_14_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_15_scaledX = {{2'd0}, ans_15[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_15_sum = io_featuresOut_15_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_15_minVal = io_featuresOut_15_sum < 8'h40 ? io_featuresOut_15_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_16_scaledX = {{2'd0}, ans_16[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_16_sum = io_featuresOut_16_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_16_minVal = io_featuresOut_16_sum < 8'h40 ? io_featuresOut_16_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_17_scaledX = {{2'd0}, ans_17[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_17_sum = io_featuresOut_17_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_17_minVal = io_featuresOut_17_sum < 8'h40 ? io_featuresOut_17_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_18_scaledX = {{2'd0}, ans_18[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_18_sum = io_featuresOut_18_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_18_minVal = io_featuresOut_18_sum < 8'h40 ? io_featuresOut_18_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_19_scaledX = {{2'd0}, ans_19[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_19_sum = io_featuresOut_19_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_19_minVal = io_featuresOut_19_sum < 8'h40 ? io_featuresOut_19_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_20_scaledX = {{2'd0}, ans_20[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_20_sum = io_featuresOut_20_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_20_minVal = io_featuresOut_20_sum < 8'h40 ? io_featuresOut_20_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_21_scaledX = {{2'd0}, ans_21[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_21_sum = io_featuresOut_21_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_21_minVal = io_featuresOut_21_sum < 8'h40 ? io_featuresOut_21_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_22_scaledX = {{2'd0}, ans_22[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_22_sum = io_featuresOut_22_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_22_minVal = io_featuresOut_22_sum < 8'h40 ? io_featuresOut_22_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_23_scaledX = {{2'd0}, ans_23[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_23_sum = io_featuresOut_23_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_23_minVal = io_featuresOut_23_sum < 8'h40 ? io_featuresOut_23_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_24_scaledX = {{2'd0}, ans_24[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_24_sum = io_featuresOut_24_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_24_minVal = io_featuresOut_24_sum < 8'h40 ? io_featuresOut_24_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_25_scaledX = {{2'd0}, ans_25[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_25_sum = io_featuresOut_25_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_25_minVal = io_featuresOut_25_sum < 8'h40 ? io_featuresOut_25_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_26_scaledX = {{2'd0}, ans_26[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_26_sum = io_featuresOut_26_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_26_minVal = io_featuresOut_26_sum < 8'h40 ? io_featuresOut_26_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_27_scaledX = {{2'd0}, ans_27[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_27_sum = io_featuresOut_27_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_27_minVal = io_featuresOut_27_sum < 8'h40 ? io_featuresOut_27_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_28_scaledX = {{2'd0}, ans_28[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_28_sum = io_featuresOut_28_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_28_minVal = io_featuresOut_28_sum < 8'h40 ? io_featuresOut_28_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_29_scaledX = {{2'd0}, ans_29[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_29_sum = io_featuresOut_29_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_29_minVal = io_featuresOut_29_sum < 8'h40 ? io_featuresOut_29_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_30_scaledX = {{2'd0}, ans_30[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_30_sum = io_featuresOut_30_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_30_minVal = io_featuresOut_30_sum < 8'h40 ? io_featuresOut_30_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_31_scaledX = {{2'd0}, ans_31[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_31_sum = io_featuresOut_31_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_31_minVal = io_featuresOut_31_sum < 8'h40 ? io_featuresOut_31_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_32_scaledX = {{2'd0}, ans_32[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_32_sum = io_featuresOut_32_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_32_minVal = io_featuresOut_32_sum < 8'h40 ? io_featuresOut_32_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_33_scaledX = {{2'd0}, ans_33[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_33_sum = io_featuresOut_33_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_33_minVal = io_featuresOut_33_sum < 8'h40 ? io_featuresOut_33_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_34_scaledX = {{2'd0}, ans_34[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_34_sum = io_featuresOut_34_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_34_minVal = io_featuresOut_34_sum < 8'h40 ? io_featuresOut_34_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_35_scaledX = {{2'd0}, ans_35[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_35_sum = io_featuresOut_35_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_35_minVal = io_featuresOut_35_sum < 8'h40 ? io_featuresOut_35_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_36_scaledX = {{2'd0}, ans_36[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_36_sum = io_featuresOut_36_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_36_minVal = io_featuresOut_36_sum < 8'h40 ? io_featuresOut_36_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_37_scaledX = {{2'd0}, ans_37[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_37_sum = io_featuresOut_37_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_37_minVal = io_featuresOut_37_sum < 8'h40 ? io_featuresOut_37_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_38_scaledX = {{2'd0}, ans_38[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_38_sum = io_featuresOut_38_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_38_minVal = io_featuresOut_38_sum < 8'h40 ? io_featuresOut_38_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_39_scaledX = {{2'd0}, ans_39[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_39_sum = io_featuresOut_39_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_39_minVal = io_featuresOut_39_sum < 8'h40 ? io_featuresOut_39_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_40_scaledX = {{2'd0}, ans_40[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_40_sum = io_featuresOut_40_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_40_minVal = io_featuresOut_40_sum < 8'h40 ? io_featuresOut_40_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_41_scaledX = {{2'd0}, ans_41[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_41_sum = io_featuresOut_41_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_41_minVal = io_featuresOut_41_sum < 8'h40 ? io_featuresOut_41_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_42_scaledX = {{2'd0}, ans_42[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_42_sum = io_featuresOut_42_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_42_minVal = io_featuresOut_42_sum < 8'h40 ? io_featuresOut_42_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_43_scaledX = {{2'd0}, ans_43[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_43_sum = io_featuresOut_43_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_43_minVal = io_featuresOut_43_sum < 8'h40 ? io_featuresOut_43_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_44_scaledX = {{2'd0}, ans_44[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_44_sum = io_featuresOut_44_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_44_minVal = io_featuresOut_44_sum < 8'h40 ? io_featuresOut_44_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_45_scaledX = {{2'd0}, ans_45[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_45_sum = io_featuresOut_45_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_45_minVal = io_featuresOut_45_sum < 8'h40 ? io_featuresOut_45_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_46_scaledX = {{2'd0}, ans_46[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_46_sum = io_featuresOut_46_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_46_minVal = io_featuresOut_46_sum < 8'h40 ? io_featuresOut_46_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_47_scaledX = {{2'd0}, ans_47[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_47_sum = io_featuresOut_47_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_47_minVal = io_featuresOut_47_sum < 8'h40 ? io_featuresOut_47_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_48_scaledX = {{2'd0}, ans_48[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_48_sum = io_featuresOut_48_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_48_minVal = io_featuresOut_48_sum < 8'h40 ? io_featuresOut_48_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_49_scaledX = {{2'd0}, ans_49[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_49_sum = io_featuresOut_49_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_49_minVal = io_featuresOut_49_sum < 8'h40 ? io_featuresOut_49_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_50_scaledX = {{2'd0}, ans_50[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_50_sum = io_featuresOut_50_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_50_minVal = io_featuresOut_50_sum < 8'h40 ? io_featuresOut_50_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_51_scaledX = {{2'd0}, ans_51[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_51_sum = io_featuresOut_51_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_51_minVal = io_featuresOut_51_sum < 8'h40 ? io_featuresOut_51_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_52_scaledX = {{2'd0}, ans_52[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_52_sum = io_featuresOut_52_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_52_minVal = io_featuresOut_52_sum < 8'h40 ? io_featuresOut_52_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_53_scaledX = {{2'd0}, ans_53[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_53_sum = io_featuresOut_53_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_53_minVal = io_featuresOut_53_sum < 8'h40 ? io_featuresOut_53_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_54_scaledX = {{2'd0}, ans_54[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_54_sum = io_featuresOut_54_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_54_minVal = io_featuresOut_54_sum < 8'h40 ? io_featuresOut_54_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_55_scaledX = {{2'd0}, ans_55[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_55_sum = io_featuresOut_55_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_55_minVal = io_featuresOut_55_sum < 8'h40 ? io_featuresOut_55_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_56_scaledX = {{2'd0}, ans_56[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_56_sum = io_featuresOut_56_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_56_minVal = io_featuresOut_56_sum < 8'h40 ? io_featuresOut_56_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_57_scaledX = {{2'd0}, ans_57[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_57_sum = io_featuresOut_57_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_57_minVal = io_featuresOut_57_sum < 8'h40 ? io_featuresOut_57_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_58_scaledX = {{2'd0}, ans_58[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_58_sum = io_featuresOut_58_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_58_minVal = io_featuresOut_58_sum < 8'h40 ? io_featuresOut_58_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_59_scaledX = {{2'd0}, ans_59[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_59_sum = io_featuresOut_59_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_59_minVal = io_featuresOut_59_sum < 8'h40 ? io_featuresOut_59_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_60_scaledX = {{2'd0}, ans_60[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_60_sum = io_featuresOut_60_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_60_minVal = io_featuresOut_60_sum < 8'h40 ? io_featuresOut_60_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_61_scaledX = {{2'd0}, ans_61[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_61_sum = io_featuresOut_61_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_61_minVal = io_featuresOut_61_sum < 8'h40 ? io_featuresOut_61_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_62_scaledX = {{2'd0}, ans_62[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_62_sum = io_featuresOut_62_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_62_minVal = io_featuresOut_62_sum < 8'h40 ? io_featuresOut_62_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  wire [7:0] io_featuresOut_63_scaledX = {{2'd0}, ans_63[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 109:27 110:17]
  wire [7:0] io_featuresOut_63_sum = io_featuresOut_63_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 112:24]
  wire [7:0] io_featuresOut_63_minVal = io_featuresOut_63_sum < 8'h40 ? io_featuresOut_63_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 114:25]
  reg  regs__0; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__1; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__2; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__3; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg [2047:0] regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  assign io_pipe_validOut = regs__3; // @[src/main/scala/fpga/Pipeline.scala 46:21]
  assign io_pipe_phvOut = regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 37:21]
  assign io_featuresOut_0 = io_featuresOut_0_minVal > 8'h0 ? io_featuresOut_0_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_1 = io_featuresOut_1_minVal > 8'h0 ? io_featuresOut_1_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_2 = io_featuresOut_2_minVal > 8'h0 ? io_featuresOut_2_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_3 = io_featuresOut_3_minVal > 8'h0 ? io_featuresOut_3_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_4 = io_featuresOut_4_minVal > 8'h0 ? io_featuresOut_4_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_5 = io_featuresOut_5_minVal > 8'h0 ? io_featuresOut_5_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_6 = io_featuresOut_6_minVal > 8'h0 ? io_featuresOut_6_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_7 = io_featuresOut_7_minVal > 8'h0 ? io_featuresOut_7_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_8 = io_featuresOut_8_minVal > 8'h0 ? io_featuresOut_8_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_9 = io_featuresOut_9_minVal > 8'h0 ? io_featuresOut_9_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_10 = io_featuresOut_10_minVal > 8'h0 ? io_featuresOut_10_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_11 = io_featuresOut_11_minVal > 8'h0 ? io_featuresOut_11_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_12 = io_featuresOut_12_minVal > 8'h0 ? io_featuresOut_12_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_13 = io_featuresOut_13_minVal > 8'h0 ? io_featuresOut_13_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_14 = io_featuresOut_14_minVal > 8'h0 ? io_featuresOut_14_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_15 = io_featuresOut_15_minVal > 8'h0 ? io_featuresOut_15_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_16 = io_featuresOut_16_minVal > 8'h0 ? io_featuresOut_16_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_17 = io_featuresOut_17_minVal > 8'h0 ? io_featuresOut_17_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_18 = io_featuresOut_18_minVal > 8'h0 ? io_featuresOut_18_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_19 = io_featuresOut_19_minVal > 8'h0 ? io_featuresOut_19_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_20 = io_featuresOut_20_minVal > 8'h0 ? io_featuresOut_20_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_21 = io_featuresOut_21_minVal > 8'h0 ? io_featuresOut_21_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_22 = io_featuresOut_22_minVal > 8'h0 ? io_featuresOut_22_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_23 = io_featuresOut_23_minVal > 8'h0 ? io_featuresOut_23_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_24 = io_featuresOut_24_minVal > 8'h0 ? io_featuresOut_24_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_25 = io_featuresOut_25_minVal > 8'h0 ? io_featuresOut_25_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_26 = io_featuresOut_26_minVal > 8'h0 ? io_featuresOut_26_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_27 = io_featuresOut_27_minVal > 8'h0 ? io_featuresOut_27_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_28 = io_featuresOut_28_minVal > 8'h0 ? io_featuresOut_28_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_29 = io_featuresOut_29_minVal > 8'h0 ? io_featuresOut_29_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_30 = io_featuresOut_30_minVal > 8'h0 ? io_featuresOut_30_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_31 = io_featuresOut_31_minVal > 8'h0 ? io_featuresOut_31_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_32 = io_featuresOut_32_minVal > 8'h0 ? io_featuresOut_32_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_33 = io_featuresOut_33_minVal > 8'h0 ? io_featuresOut_33_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_34 = io_featuresOut_34_minVal > 8'h0 ? io_featuresOut_34_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_35 = io_featuresOut_35_minVal > 8'h0 ? io_featuresOut_35_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_36 = io_featuresOut_36_minVal > 8'h0 ? io_featuresOut_36_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_37 = io_featuresOut_37_minVal > 8'h0 ? io_featuresOut_37_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_38 = io_featuresOut_38_minVal > 8'h0 ? io_featuresOut_38_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_39 = io_featuresOut_39_minVal > 8'h0 ? io_featuresOut_39_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_40 = io_featuresOut_40_minVal > 8'h0 ? io_featuresOut_40_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_41 = io_featuresOut_41_minVal > 8'h0 ? io_featuresOut_41_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_42 = io_featuresOut_42_minVal > 8'h0 ? io_featuresOut_42_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_43 = io_featuresOut_43_minVal > 8'h0 ? io_featuresOut_43_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_44 = io_featuresOut_44_minVal > 8'h0 ? io_featuresOut_44_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_45 = io_featuresOut_45_minVal > 8'h0 ? io_featuresOut_45_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_46 = io_featuresOut_46_minVal > 8'h0 ? io_featuresOut_46_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_47 = io_featuresOut_47_minVal > 8'h0 ? io_featuresOut_47_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_48 = io_featuresOut_48_minVal > 8'h0 ? io_featuresOut_48_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_49 = io_featuresOut_49_minVal > 8'h0 ? io_featuresOut_49_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_50 = io_featuresOut_50_minVal > 8'h0 ? io_featuresOut_50_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_51 = io_featuresOut_51_minVal > 8'h0 ? io_featuresOut_51_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_52 = io_featuresOut_52_minVal > 8'h0 ? io_featuresOut_52_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_53 = io_featuresOut_53_minVal > 8'h0 ? io_featuresOut_53_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_54 = io_featuresOut_54_minVal > 8'h0 ? io_featuresOut_54_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_55 = io_featuresOut_55_minVal > 8'h0 ? io_featuresOut_55_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_56 = io_featuresOut_56_minVal > 8'h0 ? io_featuresOut_56_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_57 = io_featuresOut_57_minVal > 8'h0 ? io_featuresOut_57_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_58 = io_featuresOut_58_minVal > 8'h0 ? io_featuresOut_58_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_59 = io_featuresOut_59_minVal > 8'h0 ? io_featuresOut_59_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_60 = io_featuresOut_60_minVal > 8'h0 ? io_featuresOut_60_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_61 = io_featuresOut_61_minVal > 8'h0 ? io_featuresOut_61_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_62 = io_featuresOut_62_minVal > 8'h0 ? io_featuresOut_62_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  assign io_featuresOut_63 = io_featuresOut_63_minVal > 8'h0 ? io_featuresOut_63_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 115:25]
  always @(posedge clock) begin
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h0 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_0 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_1 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_2 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_3 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h4 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_4 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h5 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_5 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h6 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_6 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h7 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_7 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h8 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_8 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h9 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_9 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'ha == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_10 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'hb == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_11 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'hc == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_12 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'hd == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_13 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'he == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_14 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'hf == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_15 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h10 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_16 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h11 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_17 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h12 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_18 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h13 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_19 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h14 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_20 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h15 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_21 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h16 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_22 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h17 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_23 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h18 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_24 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h19 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_25 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1a == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_26 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1b == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_27 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1c == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_28 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1d == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_29 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1e == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_30 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h1f == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h20 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_32 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h21 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_33 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h22 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_34 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h23 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_35 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h24 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_36 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h25 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_37 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h26 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_38 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h27 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_39 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h28 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_40 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h29 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_41 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2a == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_42 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2b == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_43 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2c == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_44 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2d == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_45 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2e == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_46 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h2f == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_47 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h30 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_48 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h31 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_49 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h32 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_50 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h33 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_51 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h34 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_52 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h35 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_53 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h36 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_54 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h37 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_55 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h38 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_56 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h39 == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_57 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3a == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_58 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3b == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_59 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3c == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_60 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3d == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_61 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3e == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_62 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (5'h1f == io_config_i[4:0] & 6'h3f == io_config_j[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
          linear_weight_31_63 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 22:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h0 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_0 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_1 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_2 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_3 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h4 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_4 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h5 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_5 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h6 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_6 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h7 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_7 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h8 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_8 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h9 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_9 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'ha == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_10 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'hb == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_11 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'hc == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_12 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'hd == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_13 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'he == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_14 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'hf == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_15 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h10 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_16 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h11 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_17 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h12 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_18 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h13 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_19 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h14 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_20 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h15 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_21 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h16 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_22 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h17 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_23 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h18 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_24 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h19 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_25 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1a == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_26 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1b == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_27 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1c == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_28 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1d == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_29 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1e == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_30 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h1f == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h20 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_32 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h21 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_33 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h22 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_34 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h23 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_35 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h24 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_36 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h25 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_37 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h26 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_38 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h27 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_39 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h28 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_40 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h29 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_41 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2a == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_42 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2b == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_43 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2c == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_44 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2d == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_45 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2e == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_46 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h2f == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_47 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h30 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_48 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h31 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_49 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h32 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_50 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h33 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_51 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h34 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_52 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h35 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_53 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h36 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_54 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h37 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_55 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h38 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_56 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h39 == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_57 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3a == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_58 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3b == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_59 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3c == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_60 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3d == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_61 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3e == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_62 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 20:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:33]
        if (6'h3f == io_config_i[5:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
          linear_bias_63 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 24:38]
        end
      end
    end
    ansAll_31_0 <= ansAll_31_0_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_1 <= ansAll_31_1_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_2 <= ansAll_31_2_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_3 <= ansAll_31_3_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_4 <= ansAll_31_4_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_5 <= ansAll_31_5_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_6 <= ansAll_31_6_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_7 <= ansAll_31_7_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_8 <= ansAll_31_8_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_9 <= ansAll_31_9_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_10 <= ansAll_31_10_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_11 <= ansAll_31_11_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_12 <= ansAll_31_12_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_13 <= ansAll_31_13_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_14 <= ansAll_31_14_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_15 <= ansAll_31_15_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_16 <= ansAll_31_16_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_17 <= ansAll_31_17_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_18 <= ansAll_31_18_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_19 <= ansAll_31_19_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_20 <= ansAll_31_20_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_21 <= ansAll_31_21_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_22 <= ansAll_31_22_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_23 <= ansAll_31_23_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_24 <= ansAll_31_24_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_25 <= ansAll_31_25_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_26 <= ansAll_31_26_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_27 <= ansAll_31_27_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_28 <= ansAll_31_28_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_29 <= ansAll_31_29_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_30 <= ansAll_31_30_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_31 <= ansAll_31_31_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_32 <= ansAll_31_32_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_33 <= ansAll_31_33_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_34 <= ansAll_31_34_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_35 <= ansAll_31_35_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_36 <= ansAll_31_36_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_37 <= ansAll_31_37_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_38 <= ansAll_31_38_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_39 <= ansAll_31_39_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_40 <= ansAll_31_40_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_41 <= ansAll_31_41_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_42 <= ansAll_31_42_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_43 <= ansAll_31_43_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_44 <= ansAll_31_44_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_45 <= ansAll_31_45_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_46 <= ansAll_31_46_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_47 <= ansAll_31_47_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_48 <= ansAll_31_48_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_49 <= ansAll_31_49_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_50 <= ansAll_31_50_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_51 <= ansAll_31_51_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_52 <= ansAll_31_52_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_53 <= ansAll_31_53_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_54 <= ansAll_31_54_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_55 <= ansAll_31_55_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_56 <= ansAll_31_56_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_57 <= ansAll_31_57_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_58 <= ansAll_31_58_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_59 <= ansAll_31_59_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_60 <= ansAll_31_60_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_61 <= ansAll_31_61_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_62 <= ansAll_31_62_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    ansAll_31_63 <= ansAll_31_63_product[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 78:26]
    if (ans_0_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_0 <= 8'h0;
    end else begin
      ans_0 <= ans_0_fp8;
    end
    if (ans_1_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_1 <= 8'h0;
    end else begin
      ans_1 <= ans_1_fp8;
    end
    if (ans_2_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_2 <= 8'h0;
    end else begin
      ans_2 <= ans_2_fp8;
    end
    if (ans_3_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_3 <= 8'h0;
    end else begin
      ans_3 <= ans_3_fp8;
    end
    if (ans_4_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_4 <= 8'h0;
    end else begin
      ans_4 <= ans_4_fp8;
    end
    if (ans_5_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_5 <= 8'h0;
    end else begin
      ans_5 <= ans_5_fp8;
    end
    if (ans_6_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_6 <= 8'h0;
    end else begin
      ans_6 <= ans_6_fp8;
    end
    if (ans_7_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_7 <= 8'h0;
    end else begin
      ans_7 <= ans_7_fp8;
    end
    if (ans_8_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_8 <= 8'h0;
    end else begin
      ans_8 <= ans_8_fp8;
    end
    if (ans_9_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_9 <= 8'h0;
    end else begin
      ans_9 <= ans_9_fp8;
    end
    if (ans_10_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_10 <= 8'h0;
    end else begin
      ans_10 <= ans_10_fp8;
    end
    if (ans_11_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_11 <= 8'h0;
    end else begin
      ans_11 <= ans_11_fp8;
    end
    if (ans_12_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_12 <= 8'h0;
    end else begin
      ans_12 <= ans_12_fp8;
    end
    if (ans_13_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_13 <= 8'h0;
    end else begin
      ans_13 <= ans_13_fp8;
    end
    if (ans_14_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_14 <= 8'h0;
    end else begin
      ans_14 <= ans_14_fp8;
    end
    if (ans_15_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_15 <= 8'h0;
    end else begin
      ans_15 <= ans_15_fp8;
    end
    if (ans_16_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_16 <= 8'h0;
    end else begin
      ans_16 <= ans_16_fp8;
    end
    if (ans_17_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_17 <= 8'h0;
    end else begin
      ans_17 <= ans_17_fp8;
    end
    if (ans_18_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_18 <= 8'h0;
    end else begin
      ans_18 <= ans_18_fp8;
    end
    if (ans_19_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_19 <= 8'h0;
    end else begin
      ans_19 <= ans_19_fp8;
    end
    if (ans_20_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_20 <= 8'h0;
    end else begin
      ans_20 <= ans_20_fp8;
    end
    if (ans_21_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_21 <= 8'h0;
    end else begin
      ans_21 <= ans_21_fp8;
    end
    if (ans_22_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_22 <= 8'h0;
    end else begin
      ans_22 <= ans_22_fp8;
    end
    if (ans_23_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_23 <= 8'h0;
    end else begin
      ans_23 <= ans_23_fp8;
    end
    if (ans_24_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_24 <= 8'h0;
    end else begin
      ans_24 <= ans_24_fp8;
    end
    if (ans_25_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_25 <= 8'h0;
    end else begin
      ans_25 <= ans_25_fp8;
    end
    if (ans_26_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_26 <= 8'h0;
    end else begin
      ans_26 <= ans_26_fp8;
    end
    if (ans_27_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_27 <= 8'h0;
    end else begin
      ans_27 <= ans_27_fp8;
    end
    if (ans_28_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_28 <= 8'h0;
    end else begin
      ans_28 <= ans_28_fp8;
    end
    if (ans_29_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_29 <= 8'h0;
    end else begin
      ans_29 <= ans_29_fp8;
    end
    if (ans_30_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_30 <= 8'h0;
    end else begin
      ans_30 <= ans_30_fp8;
    end
    if (ans_31_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_31 <= 8'h0;
    end else begin
      ans_31 <= ans_31_fp8;
    end
    if (ans_32_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_32 <= 8'h0;
    end else begin
      ans_32 <= ans_32_fp8;
    end
    if (ans_33_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_33 <= 8'h0;
    end else begin
      ans_33 <= ans_33_fp8;
    end
    if (ans_34_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_34 <= 8'h0;
    end else begin
      ans_34 <= ans_34_fp8;
    end
    if (ans_35_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_35 <= 8'h0;
    end else begin
      ans_35 <= ans_35_fp8;
    end
    if (ans_36_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_36 <= 8'h0;
    end else begin
      ans_36 <= ans_36_fp8;
    end
    if (ans_37_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_37 <= 8'h0;
    end else begin
      ans_37 <= ans_37_fp8;
    end
    if (ans_38_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_38 <= 8'h0;
    end else begin
      ans_38 <= ans_38_fp8;
    end
    if (ans_39_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_39 <= 8'h0;
    end else begin
      ans_39 <= ans_39_fp8;
    end
    if (ans_40_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_40 <= 8'h0;
    end else begin
      ans_40 <= ans_40_fp8;
    end
    if (ans_41_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_41 <= 8'h0;
    end else begin
      ans_41 <= ans_41_fp8;
    end
    if (ans_42_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_42 <= 8'h0;
    end else begin
      ans_42 <= ans_42_fp8;
    end
    if (ans_43_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_43 <= 8'h0;
    end else begin
      ans_43 <= ans_43_fp8;
    end
    if (ans_44_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_44 <= 8'h0;
    end else begin
      ans_44 <= ans_44_fp8;
    end
    if (ans_45_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_45 <= 8'h0;
    end else begin
      ans_45 <= ans_45_fp8;
    end
    if (ans_46_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_46 <= 8'h0;
    end else begin
      ans_46 <= ans_46_fp8;
    end
    if (ans_47_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_47 <= 8'h0;
    end else begin
      ans_47 <= ans_47_fp8;
    end
    if (ans_48_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_48 <= 8'h0;
    end else begin
      ans_48 <= ans_48_fp8;
    end
    if (ans_49_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_49 <= 8'h0;
    end else begin
      ans_49 <= ans_49_fp8;
    end
    if (ans_50_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_50 <= 8'h0;
    end else begin
      ans_50 <= ans_50_fp8;
    end
    if (ans_51_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_51 <= 8'h0;
    end else begin
      ans_51 <= ans_51_fp8;
    end
    if (ans_52_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_52 <= 8'h0;
    end else begin
      ans_52 <= ans_52_fp8;
    end
    if (ans_53_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_53 <= 8'h0;
    end else begin
      ans_53 <= ans_53_fp8;
    end
    if (ans_54_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_54 <= 8'h0;
    end else begin
      ans_54 <= ans_54_fp8;
    end
    if (ans_55_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_55 <= 8'h0;
    end else begin
      ans_55 <= ans_55_fp8;
    end
    if (ans_56_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_56 <= 8'h0;
    end else begin
      ans_56 <= ans_56_fp8;
    end
    if (ans_57_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_57 <= 8'h0;
    end else begin
      ans_57 <= ans_57_fp8;
    end
    if (ans_58_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_58 <= 8'h0;
    end else begin
      ans_58 <= ans_58_fp8;
    end
    if (ans_59_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_59 <= 8'h0;
    end else begin
      ans_59 <= ans_59_fp8;
    end
    if (ans_60_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_60 <= 8'h0;
    end else begin
      ans_60 <= ans_60_fp8;
    end
    if (ans_61_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_61 <= 8'h0;
    end else begin
      ans_61 <= ans_61_fp8;
    end
    if (ans_62_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_62 <= 8'h0;
    end else begin
      ans_62 <= ans_62_fp8;
    end
    if (ans_63_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 69:12]
      ans_63 <= 8'h0;
    end else begin
      ans_63 <= ans_63_fp8;
    end
    tempSum_0 <= tempSum_0 + ansAll_31_0; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_1 <= tempSum_1 + ansAll_31_1; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_2 <= tempSum_2 + ansAll_31_2; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_3 <= tempSum_3 + ansAll_31_3; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_4 <= tempSum_4 + ansAll_31_4; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_5 <= tempSum_5 + ansAll_31_5; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_6 <= tempSum_6 + ansAll_31_6; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_7 <= tempSum_7 + ansAll_31_7; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_8 <= tempSum_8 + ansAll_31_8; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_9 <= tempSum_9 + ansAll_31_9; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_10 <= tempSum_10 + ansAll_31_10; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_11 <= tempSum_11 + ansAll_31_11; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_12 <= tempSum_12 + ansAll_31_12; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_13 <= tempSum_13 + ansAll_31_13; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_14 <= tempSum_14 + ansAll_31_14; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_15 <= tempSum_15 + ansAll_31_15; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_16 <= tempSum_16 + ansAll_31_16; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_17 <= tempSum_17 + ansAll_31_17; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_18 <= tempSum_18 + ansAll_31_18; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_19 <= tempSum_19 + ansAll_31_19; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_20 <= tempSum_20 + ansAll_31_20; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_21 <= tempSum_21 + ansAll_31_21; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_22 <= tempSum_22 + ansAll_31_22; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_23 <= tempSum_23 + ansAll_31_23; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_24 <= tempSum_24 + ansAll_31_24; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_25 <= tempSum_25 + ansAll_31_25; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_26 <= tempSum_26 + ansAll_31_26; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_27 <= tempSum_27 + ansAll_31_27; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_28 <= tempSum_28 + ansAll_31_28; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_29 <= tempSum_29 + ansAll_31_29; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_30 <= tempSum_30 + ansAll_31_30; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_31 <= tempSum_31 + ansAll_31_31; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_32 <= tempSum_32 + ansAll_31_32; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_33 <= tempSum_33 + ansAll_31_33; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_34 <= tempSum_34 + ansAll_31_34; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_35 <= tempSum_35 + ansAll_31_35; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_36 <= tempSum_36 + ansAll_31_36; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_37 <= tempSum_37 + ansAll_31_37; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_38 <= tempSum_38 + ansAll_31_38; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_39 <= tempSum_39 + ansAll_31_39; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_40 <= tempSum_40 + ansAll_31_40; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_41 <= tempSum_41 + ansAll_31_41; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_42 <= tempSum_42 + ansAll_31_42; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_43 <= tempSum_43 + ansAll_31_43; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_44 <= tempSum_44 + ansAll_31_44; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_45 <= tempSum_45 + ansAll_31_45; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_46 <= tempSum_46 + ansAll_31_46; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_47 <= tempSum_47 + ansAll_31_47; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_48 <= tempSum_48 + ansAll_31_48; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_49 <= tempSum_49 + ansAll_31_49; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_50 <= tempSum_50 + ansAll_31_50; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_51 <= tempSum_51 + ansAll_31_51; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_52 <= tempSum_52 + ansAll_31_52; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_53 <= tempSum_53 + ansAll_31_53; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_54 <= tempSum_54 + ansAll_31_54; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_55 <= tempSum_55 + ansAll_31_55; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_56 <= tempSum_56 + ansAll_31_56; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_57 <= tempSum_57 + ansAll_31_57; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_58 <= tempSum_58 + ansAll_31_58; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_59 <= tempSum_59 + ansAll_31_59; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_60 <= tempSum_60 + ansAll_31_60; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_61 <= tempSum_61 + ansAll_31_61; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_62 <= tempSum_62 + ansAll_31_62; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    tempSum_63 <= tempSum_63 + ansAll_31_63; // @[src/main/scala/Multiple/LinearCompute.scala 94:38]
    regs__0 <= io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 45:25]
    regs__1 <= regs__0; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__2 <= regs__1; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__3 <= regs__2; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs_1_0 <= io_pipe_phvIn; // @[src/main/scala/fpga/Pipeline.scala 36:25]
    regs_1_1 <= regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_2 <= regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_3 <= regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 34:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  linear_weight_31_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  linear_weight_31_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  linear_weight_31_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  linear_weight_31_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  linear_weight_31_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  linear_weight_31_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  linear_weight_31_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  linear_weight_31_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  linear_weight_31_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  linear_weight_31_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  linear_weight_31_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  linear_weight_31_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  linear_weight_31_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  linear_weight_31_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  linear_weight_31_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  linear_weight_31_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  linear_weight_31_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  linear_weight_31_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  linear_weight_31_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  linear_weight_31_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  linear_weight_31_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  linear_weight_31_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  linear_weight_31_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  linear_weight_31_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  linear_weight_31_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  linear_weight_31_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  linear_weight_31_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  linear_weight_31_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  linear_weight_31_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  linear_weight_31_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  linear_weight_31_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  linear_weight_31_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  linear_weight_31_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  linear_weight_31_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  linear_weight_31_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  linear_weight_31_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  linear_weight_31_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  linear_weight_31_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  linear_weight_31_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  linear_weight_31_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  linear_weight_31_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  linear_weight_31_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  linear_weight_31_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  linear_weight_31_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  linear_weight_31_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  linear_weight_31_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  linear_weight_31_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  linear_weight_31_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  linear_weight_31_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  linear_weight_31_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  linear_weight_31_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  linear_weight_31_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  linear_weight_31_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  linear_weight_31_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  linear_weight_31_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  linear_weight_31_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  linear_weight_31_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  linear_weight_31_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  linear_weight_31_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  linear_weight_31_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  linear_weight_31_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  linear_weight_31_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  linear_weight_31_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  linear_weight_31_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  linear_bias_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  linear_bias_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  linear_bias_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  linear_bias_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  linear_bias_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  linear_bias_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  linear_bias_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  linear_bias_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  linear_bias_8 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  linear_bias_9 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  linear_bias_10 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  linear_bias_11 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  linear_bias_12 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  linear_bias_13 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  linear_bias_14 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  linear_bias_15 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  linear_bias_16 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  linear_bias_17 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  linear_bias_18 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  linear_bias_19 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  linear_bias_20 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  linear_bias_21 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  linear_bias_22 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  linear_bias_23 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  linear_bias_24 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  linear_bias_25 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  linear_bias_26 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  linear_bias_27 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  linear_bias_28 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  linear_bias_29 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  linear_bias_30 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  linear_bias_31 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  linear_bias_32 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  linear_bias_33 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  linear_bias_34 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  linear_bias_35 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  linear_bias_36 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  linear_bias_37 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  linear_bias_38 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  linear_bias_39 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  linear_bias_40 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  linear_bias_41 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  linear_bias_42 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  linear_bias_43 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  linear_bias_44 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  linear_bias_45 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  linear_bias_46 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  linear_bias_47 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  linear_bias_48 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  linear_bias_49 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  linear_bias_50 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  linear_bias_51 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  linear_bias_52 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  linear_bias_53 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  linear_bias_54 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  linear_bias_55 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  linear_bias_56 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  linear_bias_57 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  linear_bias_58 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  linear_bias_59 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  linear_bias_60 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  linear_bias_61 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  linear_bias_62 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  linear_bias_63 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  ansAll_31_0 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  ansAll_31_1 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  ansAll_31_2 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  ansAll_31_3 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  ansAll_31_4 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  ansAll_31_5 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  ansAll_31_6 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  ansAll_31_7 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  ansAll_31_8 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  ansAll_31_9 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  ansAll_31_10 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  ansAll_31_11 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  ansAll_31_12 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  ansAll_31_13 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  ansAll_31_14 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  ansAll_31_15 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  ansAll_31_16 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  ansAll_31_17 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  ansAll_31_18 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  ansAll_31_19 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  ansAll_31_20 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  ansAll_31_21 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  ansAll_31_22 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  ansAll_31_23 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  ansAll_31_24 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  ansAll_31_25 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  ansAll_31_26 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  ansAll_31_27 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  ansAll_31_28 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  ansAll_31_29 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  ansAll_31_30 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  ansAll_31_31 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  ansAll_31_32 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  ansAll_31_33 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  ansAll_31_34 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  ansAll_31_35 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  ansAll_31_36 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ansAll_31_37 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ansAll_31_38 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ansAll_31_39 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ansAll_31_40 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ansAll_31_41 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ansAll_31_42 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ansAll_31_43 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ansAll_31_44 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ansAll_31_45 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ansAll_31_46 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ansAll_31_47 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ansAll_31_48 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ansAll_31_49 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ansAll_31_50 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ansAll_31_51 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ansAll_31_52 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ansAll_31_53 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  ansAll_31_54 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  ansAll_31_55 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  ansAll_31_56 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  ansAll_31_57 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  ansAll_31_58 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  ansAll_31_59 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  ansAll_31_60 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  ansAll_31_61 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  ansAll_31_62 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  ansAll_31_63 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  ans_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  ans_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  ans_2 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  ans_3 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  ans_4 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  ans_5 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  ans_6 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  ans_7 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  ans_8 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  ans_9 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  ans_10 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  ans_11 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  ans_12 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  ans_13 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  ans_14 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  ans_15 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  ans_16 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  ans_17 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  ans_18 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  ans_19 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  ans_20 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  ans_21 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  ans_22 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  ans_23 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  ans_24 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  ans_25 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  ans_26 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  ans_27 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  ans_28 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  ans_29 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  ans_30 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  ans_31 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  ans_32 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  ans_33 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  ans_34 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  ans_35 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  ans_36 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  ans_37 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  ans_38 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  ans_39 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  ans_40 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  ans_41 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  ans_42 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  ans_43 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  ans_44 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  ans_45 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  ans_46 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  ans_47 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  ans_48 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  ans_49 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  ans_50 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  ans_51 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  ans_52 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  ans_53 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  ans_54 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  ans_55 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  ans_56 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  ans_57 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  ans_58 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  ans_59 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  ans_60 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  ans_61 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  ans_62 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  ans_63 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  tempSum_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  tempSum_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  tempSum_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  tempSum_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  tempSum_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  tempSum_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  tempSum_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  tempSum_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  tempSum_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  tempSum_9 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  tempSum_10 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  tempSum_11 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  tempSum_12 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  tempSum_13 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  tempSum_14 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  tempSum_15 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  tempSum_16 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  tempSum_17 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  tempSum_18 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  tempSum_19 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  tempSum_20 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  tempSum_21 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  tempSum_22 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  tempSum_23 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  tempSum_24 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  tempSum_25 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  tempSum_26 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  tempSum_27 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  tempSum_28 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  tempSum_29 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  tempSum_30 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  tempSum_31 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  tempSum_32 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  tempSum_33 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  tempSum_34 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  tempSum_35 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  tempSum_36 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  tempSum_37 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  tempSum_38 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  tempSum_39 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  tempSum_40 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  tempSum_41 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  tempSum_42 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  tempSum_43 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  tempSum_44 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  tempSum_45 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  tempSum_46 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  tempSum_47 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  tempSum_48 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  tempSum_49 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  tempSum_50 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  tempSum_51 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  tempSum_52 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  tempSum_53 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  tempSum_54 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  tempSum_55 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  tempSum_56 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  tempSum_57 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  tempSum_58 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  tempSum_59 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  tempSum_60 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  tempSum_61 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  tempSum_62 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  tempSum_63 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  regs__0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  regs__1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  regs__2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  regs__3 = _RAND_323[0:0];
  _RAND_324 = {64{`RANDOM}};
  regs_1_0 = _RAND_324[2047:0];
  _RAND_325 = {64{`RANDOM}};
  regs_1_1 = _RAND_325[2047:0];
  _RAND_326 = {64{`RANDOM}};
  regs_1_2 = _RAND_326[2047:0];
  _RAND_327 = {64{`RANDOM}};
  regs_1_3 = _RAND_327[2047:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAELoss(
  input           clock,
  input  [7:0]    io_featuresIn_0, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_1, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_2, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_3, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_4, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_5, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_6, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_7, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_8, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_9, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_10, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_11, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_12, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_13, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_14, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_15, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_16, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_17, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_18, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_19, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_20, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_21, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_22, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_23, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_24, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_25, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_26, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_27, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_28, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_29, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_30, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_31, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_32, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_33, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_34, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_35, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_36, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_37, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_38, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_39, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_40, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_41, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_42, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_43, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_44, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_45, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_46, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_47, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_48, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_49, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_50, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_51, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_52, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_53, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_54, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_55, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_56, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_57, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_58, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_59, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_60, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_61, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_62, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [7:0]    io_featuresIn_63, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input           io_pipe_validIn, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  output          io_pipe_validOut, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/fpga/MAELoss.scala 6:20]
  output [15:0]   io_ans // @[src/main/scala/fpga/MAELoss.scala 6:20]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [2047:0] _RAND_76;
  reg [2047:0] _RAND_77;
  reg [2047:0] _RAND_78;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] mae_0; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_1; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_2; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_3; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_4; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_5; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_6; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_7; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_8; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_9; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_10; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_11; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_12; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_13; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_14; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_15; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_16; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_17; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_18; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_19; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_20; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_21; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_22; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_23; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_24; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_25; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_26; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_27; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_28; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_29; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_30; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_31; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_32; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_33; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_34; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_35; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_36; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_37; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_38; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_39; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_40; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_41; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_42; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_43; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_44; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_45; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_46; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_47; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_48; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_49; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_50; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_51; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_52; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_53; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_54; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_55; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_56; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_57; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_58; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_59; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_60; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_61; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_62; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  reg [15:0] mae_63; // @[src/main/scala/fpga/MAELoss.scala 12:22]
  wire [7:0] featuresOriginal_0 = io_pipe_phvIn[343:336]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_1 = io_pipe_phvIn[351:344]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_2 = io_pipe_phvIn[359:352]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_3 = io_pipe_phvIn[367:360]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_4 = io_pipe_phvIn[375:368]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_5 = io_pipe_phvIn[383:376]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_6 = io_pipe_phvIn[391:384]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_7 = io_pipe_phvIn[399:392]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_8 = io_pipe_phvIn[407:400]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_9 = io_pipe_phvIn[415:408]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_10 = io_pipe_phvIn[423:416]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_11 = io_pipe_phvIn[431:424]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_12 = io_pipe_phvIn[439:432]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_13 = io_pipe_phvIn[447:440]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_14 = io_pipe_phvIn[455:448]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_15 = io_pipe_phvIn[463:456]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_16 = io_pipe_phvIn[471:464]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_17 = io_pipe_phvIn[479:472]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_18 = io_pipe_phvIn[487:480]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_19 = io_pipe_phvIn[495:488]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_20 = io_pipe_phvIn[503:496]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_21 = io_pipe_phvIn[511:504]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_22 = io_pipe_phvIn[519:512]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_23 = io_pipe_phvIn[527:520]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_24 = io_pipe_phvIn[535:528]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_25 = io_pipe_phvIn[543:536]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_26 = io_pipe_phvIn[551:544]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_27 = io_pipe_phvIn[559:552]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_28 = io_pipe_phvIn[567:560]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_29 = io_pipe_phvIn[575:568]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_30 = io_pipe_phvIn[583:576]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_31 = io_pipe_phvIn[591:584]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_32 = io_pipe_phvIn[599:592]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_33 = io_pipe_phvIn[607:600]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_34 = io_pipe_phvIn[615:608]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_35 = io_pipe_phvIn[623:616]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_36 = io_pipe_phvIn[631:624]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_37 = io_pipe_phvIn[639:632]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_38 = io_pipe_phvIn[647:640]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_39 = io_pipe_phvIn[655:648]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_40 = io_pipe_phvIn[663:656]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_41 = io_pipe_phvIn[671:664]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_42 = io_pipe_phvIn[679:672]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_43 = io_pipe_phvIn[687:680]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_44 = io_pipe_phvIn[695:688]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_45 = io_pipe_phvIn[703:696]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_46 = io_pipe_phvIn[711:704]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_47 = io_pipe_phvIn[719:712]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_48 = io_pipe_phvIn[727:720]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_49 = io_pipe_phvIn[735:728]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_50 = io_pipe_phvIn[743:736]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_51 = io_pipe_phvIn[751:744]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_52 = io_pipe_phvIn[759:752]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_53 = io_pipe_phvIn[767:760]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_54 = io_pipe_phvIn[775:768]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_55 = io_pipe_phvIn[783:776]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_56 = io_pipe_phvIn[791:784]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_57 = io_pipe_phvIn[799:792]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_58 = io_pipe_phvIn[807:800]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_59 = io_pipe_phvIn[815:808]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_60 = io_pipe_phvIn[823:816]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_61 = io_pipe_phvIn[831:824]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_62 = io_pipe_phvIn[839:832]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] featuresOriginal_63 = io_pipe_phvIn[847:840]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  wire [7:0] _mae_0_T_1 = io_featuresIn_0 - featuresOriginal_0; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_0_T_3 = featuresOriginal_0 - io_featuresIn_0; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_0 = io_featuresIn_0 > featuresOriginal_0 ? _mae_0_T_1 : _mae_0_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_1_T_1 = io_featuresIn_1 - featuresOriginal_1; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_1_T_3 = featuresOriginal_1 - io_featuresIn_1; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_1 = io_featuresIn_1 > featuresOriginal_1 ? _mae_1_T_1 : _mae_1_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_2_T_1 = io_featuresIn_2 - featuresOriginal_2; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_2_T_3 = featuresOriginal_2 - io_featuresIn_2; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_2 = io_featuresIn_2 > featuresOriginal_2 ? _mae_2_T_1 : _mae_2_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_3_T_1 = io_featuresIn_3 - featuresOriginal_3; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_3_T_3 = featuresOriginal_3 - io_featuresIn_3; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_3 = io_featuresIn_3 > featuresOriginal_3 ? _mae_3_T_1 : _mae_3_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_4_T_1 = io_featuresIn_4 - featuresOriginal_4; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_4_T_3 = featuresOriginal_4 - io_featuresIn_4; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_4 = io_featuresIn_4 > featuresOriginal_4 ? _mae_4_T_1 : _mae_4_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_5_T_1 = io_featuresIn_5 - featuresOriginal_5; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_5_T_3 = featuresOriginal_5 - io_featuresIn_5; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_5 = io_featuresIn_5 > featuresOriginal_5 ? _mae_5_T_1 : _mae_5_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_6_T_1 = io_featuresIn_6 - featuresOriginal_6; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_6_T_3 = featuresOriginal_6 - io_featuresIn_6; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_6 = io_featuresIn_6 > featuresOriginal_6 ? _mae_6_T_1 : _mae_6_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_7_T_1 = io_featuresIn_7 - featuresOriginal_7; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_7_T_3 = featuresOriginal_7 - io_featuresIn_7; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_7 = io_featuresIn_7 > featuresOriginal_7 ? _mae_7_T_1 : _mae_7_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_8_T_1 = io_featuresIn_8 - featuresOriginal_8; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_8_T_3 = featuresOriginal_8 - io_featuresIn_8; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_8 = io_featuresIn_8 > featuresOriginal_8 ? _mae_8_T_1 : _mae_8_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_9_T_1 = io_featuresIn_9 - featuresOriginal_9; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_9_T_3 = featuresOriginal_9 - io_featuresIn_9; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_9 = io_featuresIn_9 > featuresOriginal_9 ? _mae_9_T_1 : _mae_9_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_10_T_1 = io_featuresIn_10 - featuresOriginal_10; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_10_T_3 = featuresOriginal_10 - io_featuresIn_10; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_10 = io_featuresIn_10 > featuresOriginal_10 ? _mae_10_T_1 : _mae_10_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_11_T_1 = io_featuresIn_11 - featuresOriginal_11; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_11_T_3 = featuresOriginal_11 - io_featuresIn_11; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_11 = io_featuresIn_11 > featuresOriginal_11 ? _mae_11_T_1 : _mae_11_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_12_T_1 = io_featuresIn_12 - featuresOriginal_12; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_12_T_3 = featuresOriginal_12 - io_featuresIn_12; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_12 = io_featuresIn_12 > featuresOriginal_12 ? _mae_12_T_1 : _mae_12_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_13_T_1 = io_featuresIn_13 - featuresOriginal_13; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_13_T_3 = featuresOriginal_13 - io_featuresIn_13; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_13 = io_featuresIn_13 > featuresOriginal_13 ? _mae_13_T_1 : _mae_13_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_14_T_1 = io_featuresIn_14 - featuresOriginal_14; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_14_T_3 = featuresOriginal_14 - io_featuresIn_14; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_14 = io_featuresIn_14 > featuresOriginal_14 ? _mae_14_T_1 : _mae_14_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_15_T_1 = io_featuresIn_15 - featuresOriginal_15; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_15_T_3 = featuresOriginal_15 - io_featuresIn_15; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_15 = io_featuresIn_15 > featuresOriginal_15 ? _mae_15_T_1 : _mae_15_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_16_T_1 = io_featuresIn_16 - featuresOriginal_16; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_16_T_3 = featuresOriginal_16 - io_featuresIn_16; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_16 = io_featuresIn_16 > featuresOriginal_16 ? _mae_16_T_1 : _mae_16_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_17_T_1 = io_featuresIn_17 - featuresOriginal_17; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_17_T_3 = featuresOriginal_17 - io_featuresIn_17; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_17 = io_featuresIn_17 > featuresOriginal_17 ? _mae_17_T_1 : _mae_17_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_18_T_1 = io_featuresIn_18 - featuresOriginal_18; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_18_T_3 = featuresOriginal_18 - io_featuresIn_18; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_18 = io_featuresIn_18 > featuresOriginal_18 ? _mae_18_T_1 : _mae_18_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_19_T_1 = io_featuresIn_19 - featuresOriginal_19; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_19_T_3 = featuresOriginal_19 - io_featuresIn_19; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_19 = io_featuresIn_19 > featuresOriginal_19 ? _mae_19_T_1 : _mae_19_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_20_T_1 = io_featuresIn_20 - featuresOriginal_20; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_20_T_3 = featuresOriginal_20 - io_featuresIn_20; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_20 = io_featuresIn_20 > featuresOriginal_20 ? _mae_20_T_1 : _mae_20_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_21_T_1 = io_featuresIn_21 - featuresOriginal_21; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_21_T_3 = featuresOriginal_21 - io_featuresIn_21; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_21 = io_featuresIn_21 > featuresOriginal_21 ? _mae_21_T_1 : _mae_21_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_22_T_1 = io_featuresIn_22 - featuresOriginal_22; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_22_T_3 = featuresOriginal_22 - io_featuresIn_22; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_22 = io_featuresIn_22 > featuresOriginal_22 ? _mae_22_T_1 : _mae_22_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_23_T_1 = io_featuresIn_23 - featuresOriginal_23; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_23_T_3 = featuresOriginal_23 - io_featuresIn_23; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_23 = io_featuresIn_23 > featuresOriginal_23 ? _mae_23_T_1 : _mae_23_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_24_T_1 = io_featuresIn_24 - featuresOriginal_24; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_24_T_3 = featuresOriginal_24 - io_featuresIn_24; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_24 = io_featuresIn_24 > featuresOriginal_24 ? _mae_24_T_1 : _mae_24_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_25_T_1 = io_featuresIn_25 - featuresOriginal_25; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_25_T_3 = featuresOriginal_25 - io_featuresIn_25; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_25 = io_featuresIn_25 > featuresOriginal_25 ? _mae_25_T_1 : _mae_25_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_26_T_1 = io_featuresIn_26 - featuresOriginal_26; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_26_T_3 = featuresOriginal_26 - io_featuresIn_26; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_26 = io_featuresIn_26 > featuresOriginal_26 ? _mae_26_T_1 : _mae_26_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_27_T_1 = io_featuresIn_27 - featuresOriginal_27; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_27_T_3 = featuresOriginal_27 - io_featuresIn_27; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_27 = io_featuresIn_27 > featuresOriginal_27 ? _mae_27_T_1 : _mae_27_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_28_T_1 = io_featuresIn_28 - featuresOriginal_28; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_28_T_3 = featuresOriginal_28 - io_featuresIn_28; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_28 = io_featuresIn_28 > featuresOriginal_28 ? _mae_28_T_1 : _mae_28_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_29_T_1 = io_featuresIn_29 - featuresOriginal_29; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_29_T_3 = featuresOriginal_29 - io_featuresIn_29; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_29 = io_featuresIn_29 > featuresOriginal_29 ? _mae_29_T_1 : _mae_29_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_30_T_1 = io_featuresIn_30 - featuresOriginal_30; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_30_T_3 = featuresOriginal_30 - io_featuresIn_30; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_30 = io_featuresIn_30 > featuresOriginal_30 ? _mae_30_T_1 : _mae_30_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_31_T_1 = io_featuresIn_31 - featuresOriginal_31; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_31_T_3 = featuresOriginal_31 - io_featuresIn_31; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_31 = io_featuresIn_31 > featuresOriginal_31 ? _mae_31_T_1 : _mae_31_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_32_T_1 = io_featuresIn_32 - featuresOriginal_32; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_32_T_3 = featuresOriginal_32 - io_featuresIn_32; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_32 = io_featuresIn_32 > featuresOriginal_32 ? _mae_32_T_1 : _mae_32_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_33_T_1 = io_featuresIn_33 - featuresOriginal_33; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_33_T_3 = featuresOriginal_33 - io_featuresIn_33; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_33 = io_featuresIn_33 > featuresOriginal_33 ? _mae_33_T_1 : _mae_33_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_34_T_1 = io_featuresIn_34 - featuresOriginal_34; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_34_T_3 = featuresOriginal_34 - io_featuresIn_34; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_34 = io_featuresIn_34 > featuresOriginal_34 ? _mae_34_T_1 : _mae_34_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_35_T_1 = io_featuresIn_35 - featuresOriginal_35; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_35_T_3 = featuresOriginal_35 - io_featuresIn_35; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_35 = io_featuresIn_35 > featuresOriginal_35 ? _mae_35_T_1 : _mae_35_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_36_T_1 = io_featuresIn_36 - featuresOriginal_36; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_36_T_3 = featuresOriginal_36 - io_featuresIn_36; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_36 = io_featuresIn_36 > featuresOriginal_36 ? _mae_36_T_1 : _mae_36_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_37_T_1 = io_featuresIn_37 - featuresOriginal_37; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_37_T_3 = featuresOriginal_37 - io_featuresIn_37; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_37 = io_featuresIn_37 > featuresOriginal_37 ? _mae_37_T_1 : _mae_37_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_38_T_1 = io_featuresIn_38 - featuresOriginal_38; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_38_T_3 = featuresOriginal_38 - io_featuresIn_38; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_38 = io_featuresIn_38 > featuresOriginal_38 ? _mae_38_T_1 : _mae_38_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_39_T_1 = io_featuresIn_39 - featuresOriginal_39; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_39_T_3 = featuresOriginal_39 - io_featuresIn_39; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_39 = io_featuresIn_39 > featuresOriginal_39 ? _mae_39_T_1 : _mae_39_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_40_T_1 = io_featuresIn_40 - featuresOriginal_40; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_40_T_3 = featuresOriginal_40 - io_featuresIn_40; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_40 = io_featuresIn_40 > featuresOriginal_40 ? _mae_40_T_1 : _mae_40_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_41_T_1 = io_featuresIn_41 - featuresOriginal_41; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_41_T_3 = featuresOriginal_41 - io_featuresIn_41; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_41 = io_featuresIn_41 > featuresOriginal_41 ? _mae_41_T_1 : _mae_41_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_42_T_1 = io_featuresIn_42 - featuresOriginal_42; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_42_T_3 = featuresOriginal_42 - io_featuresIn_42; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_42 = io_featuresIn_42 > featuresOriginal_42 ? _mae_42_T_1 : _mae_42_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_43_T_1 = io_featuresIn_43 - featuresOriginal_43; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_43_T_3 = featuresOriginal_43 - io_featuresIn_43; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_43 = io_featuresIn_43 > featuresOriginal_43 ? _mae_43_T_1 : _mae_43_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_44_T_1 = io_featuresIn_44 - featuresOriginal_44; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_44_T_3 = featuresOriginal_44 - io_featuresIn_44; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_44 = io_featuresIn_44 > featuresOriginal_44 ? _mae_44_T_1 : _mae_44_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_45_T_1 = io_featuresIn_45 - featuresOriginal_45; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_45_T_3 = featuresOriginal_45 - io_featuresIn_45; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_45 = io_featuresIn_45 > featuresOriginal_45 ? _mae_45_T_1 : _mae_45_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_46_T_1 = io_featuresIn_46 - featuresOriginal_46; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_46_T_3 = featuresOriginal_46 - io_featuresIn_46; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_46 = io_featuresIn_46 > featuresOriginal_46 ? _mae_46_T_1 : _mae_46_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_47_T_1 = io_featuresIn_47 - featuresOriginal_47; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_47_T_3 = featuresOriginal_47 - io_featuresIn_47; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_47 = io_featuresIn_47 > featuresOriginal_47 ? _mae_47_T_1 : _mae_47_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_48_T_1 = io_featuresIn_48 - featuresOriginal_48; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_48_T_3 = featuresOriginal_48 - io_featuresIn_48; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_48 = io_featuresIn_48 > featuresOriginal_48 ? _mae_48_T_1 : _mae_48_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_49_T_1 = io_featuresIn_49 - featuresOriginal_49; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_49_T_3 = featuresOriginal_49 - io_featuresIn_49; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_49 = io_featuresIn_49 > featuresOriginal_49 ? _mae_49_T_1 : _mae_49_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_50_T_1 = io_featuresIn_50 - featuresOriginal_50; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_50_T_3 = featuresOriginal_50 - io_featuresIn_50; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_50 = io_featuresIn_50 > featuresOriginal_50 ? _mae_50_T_1 : _mae_50_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_51_T_1 = io_featuresIn_51 - featuresOriginal_51; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_51_T_3 = featuresOriginal_51 - io_featuresIn_51; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_51 = io_featuresIn_51 > featuresOriginal_51 ? _mae_51_T_1 : _mae_51_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_52_T_1 = io_featuresIn_52 - featuresOriginal_52; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_52_T_3 = featuresOriginal_52 - io_featuresIn_52; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_52 = io_featuresIn_52 > featuresOriginal_52 ? _mae_52_T_1 : _mae_52_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_53_T_1 = io_featuresIn_53 - featuresOriginal_53; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_53_T_3 = featuresOriginal_53 - io_featuresIn_53; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_53 = io_featuresIn_53 > featuresOriginal_53 ? _mae_53_T_1 : _mae_53_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_54_T_1 = io_featuresIn_54 - featuresOriginal_54; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_54_T_3 = featuresOriginal_54 - io_featuresIn_54; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_54 = io_featuresIn_54 > featuresOriginal_54 ? _mae_54_T_1 : _mae_54_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_55_T_1 = io_featuresIn_55 - featuresOriginal_55; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_55_T_3 = featuresOriginal_55 - io_featuresIn_55; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_55 = io_featuresIn_55 > featuresOriginal_55 ? _mae_55_T_1 : _mae_55_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_56_T_1 = io_featuresIn_56 - featuresOriginal_56; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_56_T_3 = featuresOriginal_56 - io_featuresIn_56; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_56 = io_featuresIn_56 > featuresOriginal_56 ? _mae_56_T_1 : _mae_56_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_57_T_1 = io_featuresIn_57 - featuresOriginal_57; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_57_T_3 = featuresOriginal_57 - io_featuresIn_57; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_57 = io_featuresIn_57 > featuresOriginal_57 ? _mae_57_T_1 : _mae_57_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_58_T_1 = io_featuresIn_58 - featuresOriginal_58; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_58_T_3 = featuresOriginal_58 - io_featuresIn_58; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_58 = io_featuresIn_58 > featuresOriginal_58 ? _mae_58_T_1 : _mae_58_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_59_T_1 = io_featuresIn_59 - featuresOriginal_59; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_59_T_3 = featuresOriginal_59 - io_featuresIn_59; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_59 = io_featuresIn_59 > featuresOriginal_59 ? _mae_59_T_1 : _mae_59_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_60_T_1 = io_featuresIn_60 - featuresOriginal_60; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_60_T_3 = featuresOriginal_60 - io_featuresIn_60; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_60 = io_featuresIn_60 > featuresOriginal_60 ? _mae_60_T_1 : _mae_60_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_61_T_1 = io_featuresIn_61 - featuresOriginal_61; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_61_T_3 = featuresOriginal_61 - io_featuresIn_61; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_61 = io_featuresIn_61 > featuresOriginal_61 ? _mae_61_T_1 : _mae_61_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_62_T_1 = io_featuresIn_62 - featuresOriginal_62; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_62_T_3 = featuresOriginal_62 - io_featuresIn_62; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_62 = io_featuresIn_62 > featuresOriginal_62 ? _mae_62_T_1 : _mae_62_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  wire [7:0] _mae_63_T_1 = io_featuresIn_63 - featuresOriginal_63; // @[src/main/scala/fpga/MAELoss.scala 16:52]
  wire [7:0] _mae_63_T_3 = featuresOriginal_63 - io_featuresIn_63; // @[src/main/scala/fpga/MAELoss.scala 18:55]
  wire [7:0] _GEN_63 = io_featuresIn_63 > featuresOriginal_63 ? _mae_63_T_1 : _mae_63_T_3; // @[src/main/scala/fpga/MAELoss.scala 15:63 16:32 18:32]
  reg [15:0] ans1_newAns_0; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_1; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_2; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_3; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_4; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_5; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_6; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  reg [15:0] ans1_newAns_7; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  wire [15:0] _ans1_newAns_ansWire_0_T_1 = mae_0 + mae_1; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_3 = _ans1_newAns_ansWire_0_T_1 + mae_2; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_5 = _ans1_newAns_ansWire_0_T_3 + mae_3; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_7 = _ans1_newAns_ansWire_0_T_5 + mae_4; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_9 = _ans1_newAns_ansWire_0_T_7 + mae_5; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_11 = _ans1_newAns_ansWire_0_T_9 + mae_6; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_1 = mae_8 + mae_9; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_3 = _ans1_newAns_ansWire_1_T_1 + mae_10; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_5 = _ans1_newAns_ansWire_1_T_3 + mae_11; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_7 = _ans1_newAns_ansWire_1_T_5 + mae_12; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_9 = _ans1_newAns_ansWire_1_T_7 + mae_13; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_1_T_11 = _ans1_newAns_ansWire_1_T_9 + mae_14; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_1 = mae_16 + mae_17; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_3 = _ans1_newAns_ansWire_2_T_1 + mae_18; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_5 = _ans1_newAns_ansWire_2_T_3 + mae_19; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_7 = _ans1_newAns_ansWire_2_T_5 + mae_20; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_9 = _ans1_newAns_ansWire_2_T_7 + mae_21; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_2_T_11 = _ans1_newAns_ansWire_2_T_9 + mae_22; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_1 = mae_24 + mae_25; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_3 = _ans1_newAns_ansWire_3_T_1 + mae_26; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_5 = _ans1_newAns_ansWire_3_T_3 + mae_27; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_7 = _ans1_newAns_ansWire_3_T_5 + mae_28; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_9 = _ans1_newAns_ansWire_3_T_7 + mae_29; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_3_T_11 = _ans1_newAns_ansWire_3_T_9 + mae_30; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_1 = mae_32 + mae_33; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_3 = _ans1_newAns_ansWire_4_T_1 + mae_34; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_5 = _ans1_newAns_ansWire_4_T_3 + mae_35; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_7 = _ans1_newAns_ansWire_4_T_5 + mae_36; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_9 = _ans1_newAns_ansWire_4_T_7 + mae_37; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_4_T_11 = _ans1_newAns_ansWire_4_T_9 + mae_38; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_1 = mae_40 + mae_41; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_3 = _ans1_newAns_ansWire_5_T_1 + mae_42; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_5 = _ans1_newAns_ansWire_5_T_3 + mae_43; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_7 = _ans1_newAns_ansWire_5_T_5 + mae_44; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_9 = _ans1_newAns_ansWire_5_T_7 + mae_45; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_5_T_11 = _ans1_newAns_ansWire_5_T_9 + mae_46; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_1 = mae_48 + mae_49; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_3 = _ans1_newAns_ansWire_6_T_1 + mae_50; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_5 = _ans1_newAns_ansWire_6_T_3 + mae_51; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_7 = _ans1_newAns_ansWire_6_T_5 + mae_52; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_9 = _ans1_newAns_ansWire_6_T_7 + mae_53; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_6_T_11 = _ans1_newAns_ansWire_6_T_9 + mae_54; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_1 = mae_56 + mae_57; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_3 = _ans1_newAns_ansWire_7_T_1 + mae_58; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_5 = _ans1_newAns_ansWire_7_T_3 + mae_59; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_7 = _ans1_newAns_ansWire_7_T_5 + mae_60; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_9 = _ans1_newAns_ansWire_7_T_7 + mae_61; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_7_T_11 = _ans1_newAns_ansWire_7_T_9 + mae_62; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  reg [15:0] ans1_0; // @[src/main/scala/fpga/MAELoss.scala 28:33]
  wire [15:0] _ans1_newAns_ansWire_0_T_15 = ans1_newAns_0 + ans1_newAns_1; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_17 = _ans1_newAns_ansWire_0_T_15 + ans1_newAns_2; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_19 = _ans1_newAns_ansWire_0_T_17 + ans1_newAns_3; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_21 = _ans1_newAns_ansWire_0_T_19 + ans1_newAns_4; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_23 = _ans1_newAns_ansWire_0_T_21 + ans1_newAns_5; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  wire [15:0] _ans1_newAns_ansWire_0_T_25 = _ans1_newAns_ansWire_0_T_23 + ans1_newAns_6; // @[src/main/scala/fpga/MAELoss.scala 31:95]
  reg  regs__0; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__1; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__2; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg [2047:0] regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  assign io_pipe_validOut = regs__2; // @[src/main/scala/fpga/Pipeline.scala 46:21]
  assign io_pipe_phvOut = regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 37:21]
  assign io_ans = ans1_0; // @[src/main/scala/fpga/MAELoss.scala 48:16]
  always @(posedge clock) begin
    mae_0 <= {{8'd0}, _GEN_0};
    mae_1 <= {{8'd0}, _GEN_1};
    mae_2 <= {{8'd0}, _GEN_2};
    mae_3 <= {{8'd0}, _GEN_3};
    mae_4 <= {{8'd0}, _GEN_4};
    mae_5 <= {{8'd0}, _GEN_5};
    mae_6 <= {{8'd0}, _GEN_6};
    mae_7 <= {{8'd0}, _GEN_7};
    mae_8 <= {{8'd0}, _GEN_8};
    mae_9 <= {{8'd0}, _GEN_9};
    mae_10 <= {{8'd0}, _GEN_10};
    mae_11 <= {{8'd0}, _GEN_11};
    mae_12 <= {{8'd0}, _GEN_12};
    mae_13 <= {{8'd0}, _GEN_13};
    mae_14 <= {{8'd0}, _GEN_14};
    mae_15 <= {{8'd0}, _GEN_15};
    mae_16 <= {{8'd0}, _GEN_16};
    mae_17 <= {{8'd0}, _GEN_17};
    mae_18 <= {{8'd0}, _GEN_18};
    mae_19 <= {{8'd0}, _GEN_19};
    mae_20 <= {{8'd0}, _GEN_20};
    mae_21 <= {{8'd0}, _GEN_21};
    mae_22 <= {{8'd0}, _GEN_22};
    mae_23 <= {{8'd0}, _GEN_23};
    mae_24 <= {{8'd0}, _GEN_24};
    mae_25 <= {{8'd0}, _GEN_25};
    mae_26 <= {{8'd0}, _GEN_26};
    mae_27 <= {{8'd0}, _GEN_27};
    mae_28 <= {{8'd0}, _GEN_28};
    mae_29 <= {{8'd0}, _GEN_29};
    mae_30 <= {{8'd0}, _GEN_30};
    mae_31 <= {{8'd0}, _GEN_31};
    mae_32 <= {{8'd0}, _GEN_32};
    mae_33 <= {{8'd0}, _GEN_33};
    mae_34 <= {{8'd0}, _GEN_34};
    mae_35 <= {{8'd0}, _GEN_35};
    mae_36 <= {{8'd0}, _GEN_36};
    mae_37 <= {{8'd0}, _GEN_37};
    mae_38 <= {{8'd0}, _GEN_38};
    mae_39 <= {{8'd0}, _GEN_39};
    mae_40 <= {{8'd0}, _GEN_40};
    mae_41 <= {{8'd0}, _GEN_41};
    mae_42 <= {{8'd0}, _GEN_42};
    mae_43 <= {{8'd0}, _GEN_43};
    mae_44 <= {{8'd0}, _GEN_44};
    mae_45 <= {{8'd0}, _GEN_45};
    mae_46 <= {{8'd0}, _GEN_46};
    mae_47 <= {{8'd0}, _GEN_47};
    mae_48 <= {{8'd0}, _GEN_48};
    mae_49 <= {{8'd0}, _GEN_49};
    mae_50 <= {{8'd0}, _GEN_50};
    mae_51 <= {{8'd0}, _GEN_51};
    mae_52 <= {{8'd0}, _GEN_52};
    mae_53 <= {{8'd0}, _GEN_53};
    mae_54 <= {{8'd0}, _GEN_54};
    mae_55 <= {{8'd0}, _GEN_55};
    mae_56 <= {{8'd0}, _GEN_56};
    mae_57 <= {{8'd0}, _GEN_57};
    mae_58 <= {{8'd0}, _GEN_58};
    mae_59 <= {{8'd0}, _GEN_59};
    mae_60 <= {{8'd0}, _GEN_60};
    mae_61 <= {{8'd0}, _GEN_61};
    mae_62 <= {{8'd0}, _GEN_62};
    mae_63 <= {{8'd0}, _GEN_63};
    ans1_newAns_0 <= _ans1_newAns_ansWire_0_T_11 + mae_7; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_1 <= _ans1_newAns_ansWire_1_T_11 + mae_15; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_2 <= _ans1_newAns_ansWire_2_T_11 + mae_23; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_3 <= _ans1_newAns_ansWire_3_T_11 + mae_31; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_4 <= _ans1_newAns_ansWire_4_T_11 + mae_39; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_5 <= _ans1_newAns_ansWire_5_T_11 + mae_47; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_6 <= _ans1_newAns_ansWire_6_T_11 + mae_55; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_newAns_7 <= _ans1_newAns_ansWire_7_T_11 + mae_63; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    ans1_0 <= _ans1_newAns_ansWire_0_T_25 + ans1_newAns_7; // @[src/main/scala/fpga/MAELoss.scala 31:95]
    regs__0 <= io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 45:25]
    regs__1 <= regs__0; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__2 <= regs__1; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs_1_0 <= io_pipe_phvIn; // @[src/main/scala/fpga/Pipeline.scala 36:25]
    regs_1_1 <= regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_2 <= regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 34:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mae_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  mae_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  mae_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  mae_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  mae_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  mae_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  mae_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  mae_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  mae_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  mae_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  mae_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  mae_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  mae_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  mae_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  mae_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  mae_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  mae_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  mae_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  mae_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  mae_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  mae_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  mae_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  mae_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  mae_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  mae_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  mae_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  mae_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  mae_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  mae_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  mae_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  mae_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  mae_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  mae_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  mae_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  mae_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  mae_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  mae_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  mae_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  mae_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  mae_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  mae_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  mae_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  mae_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  mae_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  mae_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  mae_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  mae_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  mae_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  mae_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  mae_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  mae_50 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  mae_51 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  mae_52 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  mae_53 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  mae_54 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  mae_55 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  mae_56 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  mae_57 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  mae_58 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  mae_59 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  mae_60 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  mae_61 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  mae_62 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  mae_63 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  ans1_newAns_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  ans1_newAns_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  ans1_newAns_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  ans1_newAns_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  ans1_newAns_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  ans1_newAns_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  ans1_newAns_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  ans1_newAns_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  ans1_0 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  regs__0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  regs__1 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  regs__2 = _RAND_75[0:0];
  _RAND_76 = {64{`RANDOM}};
  regs_1_0 = _RAND_76[2047:0];
  _RAND_77 = {64{`RANDOM}};
  regs_1_1 = _RAND_77[2047:0];
  _RAND_78 = {64{`RANDOM}};
  regs_1_2 = _RAND_78[2047:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Rebuild(
  input           clock,
  input           io_pipe_validIn, // @[src/main/scala/Multiple/Rebuild.scala 8:20]
  output          io_pipe_validOut, // @[src/main/scala/Multiple/Rebuild.scala 8:20]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/Multiple/Rebuild.scala 8:20]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/Multiple/Rebuild.scala 8:20]
  input  [15:0]   io_ans // @[src/main/scala/Multiple/Rebuild.scala 8:20]
);
`ifdef RANDOMIZE_REG_INIT
  reg [1023:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1023:0] reg_; // @[src/main/scala/fpga/Pipeline.scala 11:30]
  reg  reg_1; // @[src/main/scala/fpga/Pipeline.scala 18:30]
  assign io_pipe_validOut = reg_1; // @[src/main/scala/fpga/Pipeline.scala 20:21]
  assign io_pipe_phvOut = {{1024'd0}, reg_}; // @[src/main/scala/fpga/Pipeline.scala 13:21]
  always @(posedge clock) begin
    reg_ <= {io_ans[13:6],io_pipe_phvIn[1015:0]}; // @[src/main/scala/Multiple/Rebuild.scala 13:22]
    reg_1 <= io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 19:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {32{`RANDOM}};
  reg_ = _RAND_0[1023:0];
  _RAND_1 = {1{`RANDOM}};
  reg_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input           clock,
  input           reset,
  input  [31:0]   io_addr, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [31:0]   io_data, // @[src/main/scala/Multiple/Top.scala 7:16]
  input           io_pipe_validIn, // @[src/main/scala/Multiple/Top.scala 7:16]
  output          io_pipe_validOut, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/Multiple/Top.scala 7:16]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [15:0]   io_encoderScale, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [15:0]   io_encoderZeroPoint, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [15:0]   io_decoderScale, // @[src/main/scala/Multiple/Top.scala 7:16]
  input  [15:0]   io_decoderZeroPoint // @[src/main/scala/Multiple/Top.scala 7:16]
);
  wire [31:0] ctrl_io_addr; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [31:0] ctrl_io_data; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire  ctrl_io_encoderLinearConfig_en; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire  ctrl_io_encoderLinearConfig_weight; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_encoderLinearConfig_i; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_encoderLinearConfig_j; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_encoderLinearConfig_value; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire  ctrl_io_decoderLinearConfig_en; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire  ctrl_io_decoderLinearConfig_weight; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_decoderLinearConfig_i; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_decoderLinearConfig_j; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire [7:0] ctrl_io_decoderLinearConfig_value; // @[src/main/scala/Multiple/Top.scala 17:22]
  wire  encoder_clock; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire  encoder_io_pipe_validIn; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire  encoder_io_pipe_validOut; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [2047:0] encoder_io_pipe_phvIn; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [2047:0] encoder_io_pipe_phvOut; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire  encoder_io_config_en; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire  encoder_io_config_weight; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [7:0] encoder_io_config_i; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [7:0] encoder_io_config_j; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [7:0] encoder_io_config_value; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [7:0] encoder_io_featuresIn_63; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [7:0] encoder_io_featuresOut_31; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [15:0] encoder_io_scale; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire [15:0] encoder_io_zeroPoint; // @[src/main/scala/Multiple/Top.scala 18:25]
  wire  decoder_clock; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire  decoder_io_pipe_validIn; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire  decoder_io_pipe_validOut; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [2047:0] decoder_io_pipe_phvIn; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [2047:0] decoder_io_pipe_phvOut; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire  decoder_io_config_en; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire  decoder_io_config_weight; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_config_i; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_config_j; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_config_value; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresIn_31; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_0; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_1; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_2; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_3; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_4; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_5; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_6; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_7; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_8; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_9; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_10; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_11; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_12; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_13; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_14; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_15; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_16; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_17; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_18; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_19; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_20; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_21; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_22; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_23; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_24; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_25; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_26; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_27; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_28; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_29; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_30; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_31; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_32; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_33; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_34; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_35; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_36; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_37; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_38; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_39; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_40; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_41; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_42; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_43; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_44; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_45; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_46; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_47; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_48; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_49; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_50; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_51; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_52; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_53; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_54; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_55; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_56; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_57; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_58; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_59; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_60; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_61; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_62; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [7:0] decoder_io_featuresOut_63; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [15:0] decoder_io_scale; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire [15:0] decoder_io_zeroPoint; // @[src/main/scala/Multiple/Top.scala 19:25]
  wire  maeLoss_clock; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_0; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_1; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_2; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_3; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_4; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_5; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_6; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_7; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_8; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_9; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_10; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_11; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_12; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_13; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_14; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_15; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_16; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_17; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_18; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_19; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_20; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_21; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_22; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_23; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_24; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_25; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_26; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_27; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_28; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_29; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_30; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_31; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_32; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_33; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_34; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_35; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_36; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_37; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_38; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_39; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_40; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_41; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_42; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_43; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_44; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_45; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_46; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_47; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_48; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_49; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_50; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_51; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_52; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_53; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_54; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_55; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_56; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_57; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_58; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_59; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_60; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_61; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_62; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [7:0] maeLoss_io_featuresIn_63; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire  maeLoss_io_pipe_validIn; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire  maeLoss_io_pipe_validOut; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [2047:0] maeLoss_io_pipe_phvIn; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [2047:0] maeLoss_io_pipe_phvOut; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire [15:0] maeLoss_io_ans; // @[src/main/scala/Multiple/Top.scala 20:25]
  wire  rebuild_clock; // @[src/main/scala/Multiple/Top.scala 21:25]
  wire  rebuild_io_pipe_validIn; // @[src/main/scala/Multiple/Top.scala 21:25]
  wire  rebuild_io_pipe_validOut; // @[src/main/scala/Multiple/Top.scala 21:25]
  wire [2047:0] rebuild_io_pipe_phvIn; // @[src/main/scala/Multiple/Top.scala 21:25]
  wire [2047:0] rebuild_io_pipe_phvOut; // @[src/main/scala/Multiple/Top.scala 21:25]
  wire [15:0] rebuild_io_ans; // @[src/main/scala/Multiple/Top.scala 21:25]
  ControlUnit ctrl ( // @[src/main/scala/Multiple/Top.scala 17:22]
    .io_addr(ctrl_io_addr),
    .io_data(ctrl_io_data),
    .io_encoderLinearConfig_en(ctrl_io_encoderLinearConfig_en),
    .io_encoderLinearConfig_weight(ctrl_io_encoderLinearConfig_weight),
    .io_encoderLinearConfig_i(ctrl_io_encoderLinearConfig_i),
    .io_encoderLinearConfig_j(ctrl_io_encoderLinearConfig_j),
    .io_encoderLinearConfig_value(ctrl_io_encoderLinearConfig_value),
    .io_decoderLinearConfig_en(ctrl_io_decoderLinearConfig_en),
    .io_decoderLinearConfig_weight(ctrl_io_decoderLinearConfig_weight),
    .io_decoderLinearConfig_i(ctrl_io_decoderLinearConfig_i),
    .io_decoderLinearConfig_j(ctrl_io_decoderLinearConfig_j),
    .io_decoderLinearConfig_value(ctrl_io_decoderLinearConfig_value)
  );
  LinearCompute encoder ( // @[src/main/scala/Multiple/Top.scala 18:25]
    .clock(encoder_clock),
    .io_pipe_validIn(encoder_io_pipe_validIn),
    .io_pipe_validOut(encoder_io_pipe_validOut),
    .io_pipe_phvIn(encoder_io_pipe_phvIn),
    .io_pipe_phvOut(encoder_io_pipe_phvOut),
    .io_config_en(encoder_io_config_en),
    .io_config_weight(encoder_io_config_weight),
    .io_config_i(encoder_io_config_i),
    .io_config_j(encoder_io_config_j),
    .io_config_value(encoder_io_config_value),
    .io_featuresIn_63(encoder_io_featuresIn_63),
    .io_featuresOut_31(encoder_io_featuresOut_31),
    .io_scale(encoder_io_scale),
    .io_zeroPoint(encoder_io_zeroPoint)
  );
  LinearCompute_1 decoder ( // @[src/main/scala/Multiple/Top.scala 19:25]
    .clock(decoder_clock),
    .io_pipe_validIn(decoder_io_pipe_validIn),
    .io_pipe_validOut(decoder_io_pipe_validOut),
    .io_pipe_phvIn(decoder_io_pipe_phvIn),
    .io_pipe_phvOut(decoder_io_pipe_phvOut),
    .io_config_en(decoder_io_config_en),
    .io_config_weight(decoder_io_config_weight),
    .io_config_i(decoder_io_config_i),
    .io_config_j(decoder_io_config_j),
    .io_config_value(decoder_io_config_value),
    .io_featuresIn_31(decoder_io_featuresIn_31),
    .io_featuresOut_0(decoder_io_featuresOut_0),
    .io_featuresOut_1(decoder_io_featuresOut_1),
    .io_featuresOut_2(decoder_io_featuresOut_2),
    .io_featuresOut_3(decoder_io_featuresOut_3),
    .io_featuresOut_4(decoder_io_featuresOut_4),
    .io_featuresOut_5(decoder_io_featuresOut_5),
    .io_featuresOut_6(decoder_io_featuresOut_6),
    .io_featuresOut_7(decoder_io_featuresOut_7),
    .io_featuresOut_8(decoder_io_featuresOut_8),
    .io_featuresOut_9(decoder_io_featuresOut_9),
    .io_featuresOut_10(decoder_io_featuresOut_10),
    .io_featuresOut_11(decoder_io_featuresOut_11),
    .io_featuresOut_12(decoder_io_featuresOut_12),
    .io_featuresOut_13(decoder_io_featuresOut_13),
    .io_featuresOut_14(decoder_io_featuresOut_14),
    .io_featuresOut_15(decoder_io_featuresOut_15),
    .io_featuresOut_16(decoder_io_featuresOut_16),
    .io_featuresOut_17(decoder_io_featuresOut_17),
    .io_featuresOut_18(decoder_io_featuresOut_18),
    .io_featuresOut_19(decoder_io_featuresOut_19),
    .io_featuresOut_20(decoder_io_featuresOut_20),
    .io_featuresOut_21(decoder_io_featuresOut_21),
    .io_featuresOut_22(decoder_io_featuresOut_22),
    .io_featuresOut_23(decoder_io_featuresOut_23),
    .io_featuresOut_24(decoder_io_featuresOut_24),
    .io_featuresOut_25(decoder_io_featuresOut_25),
    .io_featuresOut_26(decoder_io_featuresOut_26),
    .io_featuresOut_27(decoder_io_featuresOut_27),
    .io_featuresOut_28(decoder_io_featuresOut_28),
    .io_featuresOut_29(decoder_io_featuresOut_29),
    .io_featuresOut_30(decoder_io_featuresOut_30),
    .io_featuresOut_31(decoder_io_featuresOut_31),
    .io_featuresOut_32(decoder_io_featuresOut_32),
    .io_featuresOut_33(decoder_io_featuresOut_33),
    .io_featuresOut_34(decoder_io_featuresOut_34),
    .io_featuresOut_35(decoder_io_featuresOut_35),
    .io_featuresOut_36(decoder_io_featuresOut_36),
    .io_featuresOut_37(decoder_io_featuresOut_37),
    .io_featuresOut_38(decoder_io_featuresOut_38),
    .io_featuresOut_39(decoder_io_featuresOut_39),
    .io_featuresOut_40(decoder_io_featuresOut_40),
    .io_featuresOut_41(decoder_io_featuresOut_41),
    .io_featuresOut_42(decoder_io_featuresOut_42),
    .io_featuresOut_43(decoder_io_featuresOut_43),
    .io_featuresOut_44(decoder_io_featuresOut_44),
    .io_featuresOut_45(decoder_io_featuresOut_45),
    .io_featuresOut_46(decoder_io_featuresOut_46),
    .io_featuresOut_47(decoder_io_featuresOut_47),
    .io_featuresOut_48(decoder_io_featuresOut_48),
    .io_featuresOut_49(decoder_io_featuresOut_49),
    .io_featuresOut_50(decoder_io_featuresOut_50),
    .io_featuresOut_51(decoder_io_featuresOut_51),
    .io_featuresOut_52(decoder_io_featuresOut_52),
    .io_featuresOut_53(decoder_io_featuresOut_53),
    .io_featuresOut_54(decoder_io_featuresOut_54),
    .io_featuresOut_55(decoder_io_featuresOut_55),
    .io_featuresOut_56(decoder_io_featuresOut_56),
    .io_featuresOut_57(decoder_io_featuresOut_57),
    .io_featuresOut_58(decoder_io_featuresOut_58),
    .io_featuresOut_59(decoder_io_featuresOut_59),
    .io_featuresOut_60(decoder_io_featuresOut_60),
    .io_featuresOut_61(decoder_io_featuresOut_61),
    .io_featuresOut_62(decoder_io_featuresOut_62),
    .io_featuresOut_63(decoder_io_featuresOut_63),
    .io_scale(decoder_io_scale),
    .io_zeroPoint(decoder_io_zeroPoint)
  );
  MAELoss maeLoss ( // @[src/main/scala/Multiple/Top.scala 20:25]
    .clock(maeLoss_clock),
    .io_featuresIn_0(maeLoss_io_featuresIn_0),
    .io_featuresIn_1(maeLoss_io_featuresIn_1),
    .io_featuresIn_2(maeLoss_io_featuresIn_2),
    .io_featuresIn_3(maeLoss_io_featuresIn_3),
    .io_featuresIn_4(maeLoss_io_featuresIn_4),
    .io_featuresIn_5(maeLoss_io_featuresIn_5),
    .io_featuresIn_6(maeLoss_io_featuresIn_6),
    .io_featuresIn_7(maeLoss_io_featuresIn_7),
    .io_featuresIn_8(maeLoss_io_featuresIn_8),
    .io_featuresIn_9(maeLoss_io_featuresIn_9),
    .io_featuresIn_10(maeLoss_io_featuresIn_10),
    .io_featuresIn_11(maeLoss_io_featuresIn_11),
    .io_featuresIn_12(maeLoss_io_featuresIn_12),
    .io_featuresIn_13(maeLoss_io_featuresIn_13),
    .io_featuresIn_14(maeLoss_io_featuresIn_14),
    .io_featuresIn_15(maeLoss_io_featuresIn_15),
    .io_featuresIn_16(maeLoss_io_featuresIn_16),
    .io_featuresIn_17(maeLoss_io_featuresIn_17),
    .io_featuresIn_18(maeLoss_io_featuresIn_18),
    .io_featuresIn_19(maeLoss_io_featuresIn_19),
    .io_featuresIn_20(maeLoss_io_featuresIn_20),
    .io_featuresIn_21(maeLoss_io_featuresIn_21),
    .io_featuresIn_22(maeLoss_io_featuresIn_22),
    .io_featuresIn_23(maeLoss_io_featuresIn_23),
    .io_featuresIn_24(maeLoss_io_featuresIn_24),
    .io_featuresIn_25(maeLoss_io_featuresIn_25),
    .io_featuresIn_26(maeLoss_io_featuresIn_26),
    .io_featuresIn_27(maeLoss_io_featuresIn_27),
    .io_featuresIn_28(maeLoss_io_featuresIn_28),
    .io_featuresIn_29(maeLoss_io_featuresIn_29),
    .io_featuresIn_30(maeLoss_io_featuresIn_30),
    .io_featuresIn_31(maeLoss_io_featuresIn_31),
    .io_featuresIn_32(maeLoss_io_featuresIn_32),
    .io_featuresIn_33(maeLoss_io_featuresIn_33),
    .io_featuresIn_34(maeLoss_io_featuresIn_34),
    .io_featuresIn_35(maeLoss_io_featuresIn_35),
    .io_featuresIn_36(maeLoss_io_featuresIn_36),
    .io_featuresIn_37(maeLoss_io_featuresIn_37),
    .io_featuresIn_38(maeLoss_io_featuresIn_38),
    .io_featuresIn_39(maeLoss_io_featuresIn_39),
    .io_featuresIn_40(maeLoss_io_featuresIn_40),
    .io_featuresIn_41(maeLoss_io_featuresIn_41),
    .io_featuresIn_42(maeLoss_io_featuresIn_42),
    .io_featuresIn_43(maeLoss_io_featuresIn_43),
    .io_featuresIn_44(maeLoss_io_featuresIn_44),
    .io_featuresIn_45(maeLoss_io_featuresIn_45),
    .io_featuresIn_46(maeLoss_io_featuresIn_46),
    .io_featuresIn_47(maeLoss_io_featuresIn_47),
    .io_featuresIn_48(maeLoss_io_featuresIn_48),
    .io_featuresIn_49(maeLoss_io_featuresIn_49),
    .io_featuresIn_50(maeLoss_io_featuresIn_50),
    .io_featuresIn_51(maeLoss_io_featuresIn_51),
    .io_featuresIn_52(maeLoss_io_featuresIn_52),
    .io_featuresIn_53(maeLoss_io_featuresIn_53),
    .io_featuresIn_54(maeLoss_io_featuresIn_54),
    .io_featuresIn_55(maeLoss_io_featuresIn_55),
    .io_featuresIn_56(maeLoss_io_featuresIn_56),
    .io_featuresIn_57(maeLoss_io_featuresIn_57),
    .io_featuresIn_58(maeLoss_io_featuresIn_58),
    .io_featuresIn_59(maeLoss_io_featuresIn_59),
    .io_featuresIn_60(maeLoss_io_featuresIn_60),
    .io_featuresIn_61(maeLoss_io_featuresIn_61),
    .io_featuresIn_62(maeLoss_io_featuresIn_62),
    .io_featuresIn_63(maeLoss_io_featuresIn_63),
    .io_pipe_validIn(maeLoss_io_pipe_validIn),
    .io_pipe_validOut(maeLoss_io_pipe_validOut),
    .io_pipe_phvIn(maeLoss_io_pipe_phvIn),
    .io_pipe_phvOut(maeLoss_io_pipe_phvOut),
    .io_ans(maeLoss_io_ans)
  );
  Rebuild rebuild ( // @[src/main/scala/Multiple/Top.scala 21:25]
    .clock(rebuild_clock),
    .io_pipe_validIn(rebuild_io_pipe_validIn),
    .io_pipe_validOut(rebuild_io_pipe_validOut),
    .io_pipe_phvIn(rebuild_io_pipe_phvIn),
    .io_pipe_phvOut(rebuild_io_pipe_phvOut),
    .io_ans(rebuild_io_ans)
  );
  assign io_pipe_validOut = rebuild_io_pipe_validOut; // @[src/main/scala/fpga/Pipeline.scala 82:31]
  assign io_pipe_phvOut = rebuild_io_pipe_phvOut; // @[src/main/scala/fpga/Pipeline.scala 81:29]
  assign ctrl_io_addr = io_addr; // @[src/main/scala/Multiple/Top.scala 23:18]
  assign ctrl_io_data = io_data; // @[src/main/scala/Multiple/Top.scala 24:18]
  assign encoder_clock = clock;
  assign encoder_io_pipe_validIn = io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 77:30]
  assign encoder_io_pipe_phvIn = io_pipe_phvIn; // @[src/main/scala/fpga/Pipeline.scala 76:28]
  assign encoder_io_config_en = ctrl_io_encoderLinearConfig_en; // @[src/main/scala/Multiple/Top.scala 25:33]
  assign encoder_io_config_weight = ctrl_io_encoderLinearConfig_weight; // @[src/main/scala/Multiple/Top.scala 25:33]
  assign encoder_io_config_i = ctrl_io_encoderLinearConfig_i; // @[src/main/scala/Multiple/Top.scala 25:33]
  assign encoder_io_config_j = ctrl_io_encoderLinearConfig_j; // @[src/main/scala/Multiple/Top.scala 25:33]
  assign encoder_io_config_value = ctrl_io_encoderLinearConfig_value; // @[src/main/scala/Multiple/Top.scala 25:33]
  assign encoder_io_featuresIn_63 = io_pipe_phvIn[847:840]; // @[src/main/scala/fpga/Pipeline.scala 69:70]
  assign encoder_io_scale = io_encoderScale; // @[src/main/scala/Multiple/Top.scala 28:22]
  assign encoder_io_zeroPoint = io_encoderZeroPoint; // @[src/main/scala/Multiple/Top.scala 29:26]
  assign decoder_clock = clock;
  assign decoder_io_pipe_validIn = encoder_io_pipe_validOut; // @[src/main/scala/fpga/Pipeline.scala 87:30]
  assign decoder_io_pipe_phvIn = encoder_io_pipe_phvOut; // @[src/main/scala/fpga/Pipeline.scala 86:28]
  assign decoder_io_config_en = ctrl_io_decoderLinearConfig_en; // @[src/main/scala/Multiple/Top.scala 26:33]
  assign decoder_io_config_weight = ctrl_io_decoderLinearConfig_weight; // @[src/main/scala/Multiple/Top.scala 26:33]
  assign decoder_io_config_i = ctrl_io_decoderLinearConfig_i; // @[src/main/scala/Multiple/Top.scala 26:33]
  assign decoder_io_config_j = ctrl_io_decoderLinearConfig_j; // @[src/main/scala/Multiple/Top.scala 26:33]
  assign decoder_io_config_value = ctrl_io_decoderLinearConfig_value; // @[src/main/scala/Multiple/Top.scala 26:33]
  assign decoder_io_featuresIn_31 = encoder_io_featuresOut_31; // @[src/main/scala/Multiple/Top.scala 36:27]
  assign decoder_io_scale = io_decoderScale; // @[src/main/scala/Multiple/Top.scala 30:22]
  assign decoder_io_zeroPoint = io_decoderZeroPoint; // @[src/main/scala/Multiple/Top.scala 31:26]
  assign maeLoss_clock = clock;
  assign maeLoss_io_featuresIn_0 = decoder_io_featuresOut_0; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_1 = decoder_io_featuresOut_1; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_2 = decoder_io_featuresOut_2; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_3 = decoder_io_featuresOut_3; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_4 = decoder_io_featuresOut_4; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_5 = decoder_io_featuresOut_5; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_6 = decoder_io_featuresOut_6; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_7 = decoder_io_featuresOut_7; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_8 = decoder_io_featuresOut_8; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_9 = decoder_io_featuresOut_9; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_10 = decoder_io_featuresOut_10; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_11 = decoder_io_featuresOut_11; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_12 = decoder_io_featuresOut_12; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_13 = decoder_io_featuresOut_13; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_14 = decoder_io_featuresOut_14; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_15 = decoder_io_featuresOut_15; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_16 = decoder_io_featuresOut_16; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_17 = decoder_io_featuresOut_17; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_18 = decoder_io_featuresOut_18; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_19 = decoder_io_featuresOut_19; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_20 = decoder_io_featuresOut_20; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_21 = decoder_io_featuresOut_21; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_22 = decoder_io_featuresOut_22; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_23 = decoder_io_featuresOut_23; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_24 = decoder_io_featuresOut_24; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_25 = decoder_io_featuresOut_25; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_26 = decoder_io_featuresOut_26; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_27 = decoder_io_featuresOut_27; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_28 = decoder_io_featuresOut_28; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_29 = decoder_io_featuresOut_29; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_30 = decoder_io_featuresOut_30; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_31 = decoder_io_featuresOut_31; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_32 = decoder_io_featuresOut_32; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_33 = decoder_io_featuresOut_33; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_34 = decoder_io_featuresOut_34; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_35 = decoder_io_featuresOut_35; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_36 = decoder_io_featuresOut_36; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_37 = decoder_io_featuresOut_37; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_38 = decoder_io_featuresOut_38; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_39 = decoder_io_featuresOut_39; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_40 = decoder_io_featuresOut_40; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_41 = decoder_io_featuresOut_41; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_42 = decoder_io_featuresOut_42; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_43 = decoder_io_featuresOut_43; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_44 = decoder_io_featuresOut_44; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_45 = decoder_io_featuresOut_45; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_46 = decoder_io_featuresOut_46; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_47 = decoder_io_featuresOut_47; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_48 = decoder_io_featuresOut_48; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_49 = decoder_io_featuresOut_49; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_50 = decoder_io_featuresOut_50; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_51 = decoder_io_featuresOut_51; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_52 = decoder_io_featuresOut_52; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_53 = decoder_io_featuresOut_53; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_54 = decoder_io_featuresOut_54; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_55 = decoder_io_featuresOut_55; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_56 = decoder_io_featuresOut_56; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_57 = decoder_io_featuresOut_57; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_58 = decoder_io_featuresOut_58; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_59 = decoder_io_featuresOut_59; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_60 = decoder_io_featuresOut_60; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_61 = decoder_io_featuresOut_61; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_62 = decoder_io_featuresOut_62; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_featuresIn_63 = decoder_io_featuresOut_63; // @[src/main/scala/Multiple/Top.scala 39:27]
  assign maeLoss_io_pipe_validIn = decoder_io_pipe_validOut; // @[src/main/scala/fpga/Pipeline.scala 87:30]
  assign maeLoss_io_pipe_phvIn = decoder_io_pipe_phvOut; // @[src/main/scala/fpga/Pipeline.scala 86:28]
  assign rebuild_clock = clock;
  assign rebuild_io_pipe_validIn = maeLoss_io_pipe_validOut; // @[src/main/scala/fpga/Pipeline.scala 87:30]
  assign rebuild_io_pipe_phvIn = maeLoss_io_pipe_phvOut; // @[src/main/scala/fpga/Pipeline.scala 86:28]
  assign rebuild_io_ans = maeLoss_io_ans; // @[src/main/scala/Multiple/Top.scala 42:20]
endmodule
