module LinearCompute(
  input           clock,
  input           reset,
  input           io_pipe_validIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output          io_pipe_validOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [2047:0] io_pipe_phvIn, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [2047:0] io_pipe_phvOut, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_en, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input           io_config_weight, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_i, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_j, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_config_value, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_0, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_1, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_2, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_3, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_4, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_5, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_6, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_7, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_8, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_9, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_10, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_11, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_12, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_13, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_14, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_15, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_16, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_17, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_18, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_19, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_20, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_21, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_22, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_23, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_24, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_25, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_26, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_27, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_28, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_29, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_30, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_31, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_32, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_33, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_34, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_35, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_36, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_37, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_38, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_39, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_40, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_41, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_42, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_43, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_44, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_45, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_46, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_47, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_48, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_49, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_50, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_51, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_52, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_53, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_54, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_55, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_56, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_57, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_58, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_59, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_60, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_61, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_62, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [7:0]    io_featuresIn_63, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_0, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_1, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_2, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_3, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_4, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_5, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_6, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_7, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_8, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_9, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_10, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_11, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_12, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_13, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_14, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_15, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_16, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_17, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_18, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_19, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_20, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_21, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_22, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_23, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_24, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_25, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_26, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_27, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_28, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_29, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_30, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  output [7:0]    io_featuresOut_31, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_scale, // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
  input  [15:0]   io_zeroPoint // @[src/main/scala/Multiple/LinearCompute.scala 9:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [2047:0] _RAND_196;
  reg [2047:0] _RAND_197;
  reg [2047:0] _RAND_198;
  reg [2047:0] _RAND_199;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] linear_weight_63_0; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_1; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_2; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_3; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_4; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_5; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_6; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_7; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_8; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_9; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_10; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_11; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_12; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_13; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_14; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_15; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_16; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_17; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_18; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_19; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_20; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_21; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_22; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_23; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_24; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_25; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_26; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_27; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_28; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_29; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_30; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_weight_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_0; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_1; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_2; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_3; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_4; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_5; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_6; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_7; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_8; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_9; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_10; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_11; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_12; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_13; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_14; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_15; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_16; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_17; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_18; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_19; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_20; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_21; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_22; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_23; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_24; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_25; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_26; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_27; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_28; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_29; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_30; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  reg [7:0] linear_bias_31; // @[src/main/scala/Multiple/LinearCompute.scala 18:21]
  wire [31:0] _GEN_14432 = {{16'd0}, io_zeroPoint}; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _featuresInQ8_T_126 = {24'h0,io_featuresIn_63}; // @[src/main/scala/Multiple/LinearCompute.scala 114:73]
  wire  featuresInQ8_sign_63 = _featuresInQ8_T_126[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _featuresInQ8_absX_T_189 = ~_featuresInQ8_T_126; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _featuresInQ8_absX_T_191 = _featuresInQ8_absX_T_189 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] featuresInQ8_absX_63 = featuresInQ8_sign_63 ? _featuresInQ8_absX_T_191 : _featuresInQ8_T_126; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _featuresInQ8_shiftedX_T_253 = _GEN_14432 - featuresInQ8_absX_63; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _featuresInQ8_shiftedX_T_255 = featuresInQ8_absX_63 - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] featuresInQ8_shiftedX_63 = featuresInQ8_sign_63 ? _featuresInQ8_shiftedX_T_253 :
    _featuresInQ8_shiftedX_T_255; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _featuresInQ8_scaledX_T_127 = featuresInQ8_shiftedX_63 * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] featuresInQ8_scaledX_63 = _featuresInQ8_scaledX_T_127 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _featuresInQ8_clippedX_T_191 = featuresInQ8_scaledX_63 < 49'hfffffe40 ? 49'hfffffe40 :
    featuresInQ8_scaledX_63; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] featuresInQ8_clippedX_63 = featuresInQ8_scaledX_63 > 49'h1c0 ? 49'h1c0 : _featuresInQ8_clippedX_T_191; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _featuresInQ8_absClipped_T_253 = ~featuresInQ8_clippedX_63; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _featuresInQ8_absClipped_T_255 = _featuresInQ8_absClipped_T_253 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] featuresInQ8_absClipped_63 = featuresInQ8_clippedX_63[31] ? _featuresInQ8_absClipped_T_255 :
    featuresInQ8_clippedX_63; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  featuresInQ8_isZero_63 = featuresInQ8_absClipped_63 == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_15127 = {{16'd0}, featuresInQ8_absClipped_63[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11974 = _GEN_15127 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11976 = {featuresInQ8_absClipped_63[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11978 = _featuresInQ8_leadingZeros_T_11976 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11979 = _featuresInQ8_leadingZeros_T_11974 |
    _featuresInQ8_leadingZeros_T_11978; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_15128 = {{8'd0}, _featuresInQ8_leadingZeros_T_11979[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11984 = _GEN_15128 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11986 = {_featuresInQ8_leadingZeros_T_11979[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11988 = _featuresInQ8_leadingZeros_T_11986 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11989 = _featuresInQ8_leadingZeros_T_11984 |
    _featuresInQ8_leadingZeros_T_11988; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_15129 = {{4'd0}, _featuresInQ8_leadingZeros_T_11989[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11994 = _GEN_15129 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11996 = {_featuresInQ8_leadingZeros_T_11989[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11998 = _featuresInQ8_leadingZeros_T_11996 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_11999 = _featuresInQ8_leadingZeros_T_11994 |
    _featuresInQ8_leadingZeros_T_11998; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_15130 = {{2'd0}, _featuresInQ8_leadingZeros_T_11999[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12004 = _GEN_15130 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12006 = {_featuresInQ8_leadingZeros_T_11999[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12008 = _featuresInQ8_leadingZeros_T_12006 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12009 = _featuresInQ8_leadingZeros_T_12004 |
    _featuresInQ8_leadingZeros_T_12008; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_15131 = {{1'd0}, _featuresInQ8_leadingZeros_T_12009[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12014 = _GEN_15131 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12016 = {_featuresInQ8_leadingZeros_T_12009[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12018 = _featuresInQ8_leadingZeros_T_12016 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _featuresInQ8_leadingZeros_T_12019 = _featuresInQ8_leadingZeros_T_12014 |
    _featuresInQ8_leadingZeros_T_12018; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_15132 = {{8'd0}, featuresInQ8_absClipped_63[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12025 = _GEN_15132 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12027 = {featuresInQ8_absClipped_63[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12029 = _featuresInQ8_leadingZeros_T_12027 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12030 = _featuresInQ8_leadingZeros_T_12025 |
    _featuresInQ8_leadingZeros_T_12029; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_15133 = {{4'd0}, _featuresInQ8_leadingZeros_T_12030[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12035 = _GEN_15133 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12037 = {_featuresInQ8_leadingZeros_T_12030[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12039 = _featuresInQ8_leadingZeros_T_12037 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12040 = _featuresInQ8_leadingZeros_T_12035 |
    _featuresInQ8_leadingZeros_T_12039; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_15134 = {{2'd0}, _featuresInQ8_leadingZeros_T_12040[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12045 = _GEN_15134 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12047 = {_featuresInQ8_leadingZeros_T_12040[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12049 = _featuresInQ8_leadingZeros_T_12047 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12050 = _featuresInQ8_leadingZeros_T_12045 |
    _featuresInQ8_leadingZeros_T_12049; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_15135 = {{1'd0}, _featuresInQ8_leadingZeros_T_12050[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12055 = _GEN_15135 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12057 = {_featuresInQ8_leadingZeros_T_12050[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12059 = _featuresInQ8_leadingZeros_T_12057 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _featuresInQ8_leadingZeros_T_12060 = _featuresInQ8_leadingZeros_T_12055 |
    _featuresInQ8_leadingZeros_T_12059; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _featuresInQ8_leadingZeros_T_12063 = {_featuresInQ8_leadingZeros_T_12019,
    _featuresInQ8_leadingZeros_T_12060,featuresInQ8_absClipped_63[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _featuresInQ8_leadingZeros_T_12113 = _featuresInQ8_leadingZeros_T_12063[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12114 = _featuresInQ8_leadingZeros_T_12063[46] ? 6'h2e :
    _featuresInQ8_leadingZeros_T_12113; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12115 = _featuresInQ8_leadingZeros_T_12063[45] ? 6'h2d :
    _featuresInQ8_leadingZeros_T_12114; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12116 = _featuresInQ8_leadingZeros_T_12063[44] ? 6'h2c :
    _featuresInQ8_leadingZeros_T_12115; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12117 = _featuresInQ8_leadingZeros_T_12063[43] ? 6'h2b :
    _featuresInQ8_leadingZeros_T_12116; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12118 = _featuresInQ8_leadingZeros_T_12063[42] ? 6'h2a :
    _featuresInQ8_leadingZeros_T_12117; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12119 = _featuresInQ8_leadingZeros_T_12063[41] ? 6'h29 :
    _featuresInQ8_leadingZeros_T_12118; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12120 = _featuresInQ8_leadingZeros_T_12063[40] ? 6'h28 :
    _featuresInQ8_leadingZeros_T_12119; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12121 = _featuresInQ8_leadingZeros_T_12063[39] ? 6'h27 :
    _featuresInQ8_leadingZeros_T_12120; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12122 = _featuresInQ8_leadingZeros_T_12063[38] ? 6'h26 :
    _featuresInQ8_leadingZeros_T_12121; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12123 = _featuresInQ8_leadingZeros_T_12063[37] ? 6'h25 :
    _featuresInQ8_leadingZeros_T_12122; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12124 = _featuresInQ8_leadingZeros_T_12063[36] ? 6'h24 :
    _featuresInQ8_leadingZeros_T_12123; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12125 = _featuresInQ8_leadingZeros_T_12063[35] ? 6'h23 :
    _featuresInQ8_leadingZeros_T_12124; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12126 = _featuresInQ8_leadingZeros_T_12063[34] ? 6'h22 :
    _featuresInQ8_leadingZeros_T_12125; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12127 = _featuresInQ8_leadingZeros_T_12063[33] ? 6'h21 :
    _featuresInQ8_leadingZeros_T_12126; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12128 = _featuresInQ8_leadingZeros_T_12063[32] ? 6'h20 :
    _featuresInQ8_leadingZeros_T_12127; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12129 = _featuresInQ8_leadingZeros_T_12063[31] ? 6'h1f :
    _featuresInQ8_leadingZeros_T_12128; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12130 = _featuresInQ8_leadingZeros_T_12063[30] ? 6'h1e :
    _featuresInQ8_leadingZeros_T_12129; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12131 = _featuresInQ8_leadingZeros_T_12063[29] ? 6'h1d :
    _featuresInQ8_leadingZeros_T_12130; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12132 = _featuresInQ8_leadingZeros_T_12063[28] ? 6'h1c :
    _featuresInQ8_leadingZeros_T_12131; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12133 = _featuresInQ8_leadingZeros_T_12063[27] ? 6'h1b :
    _featuresInQ8_leadingZeros_T_12132; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12134 = _featuresInQ8_leadingZeros_T_12063[26] ? 6'h1a :
    _featuresInQ8_leadingZeros_T_12133; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12135 = _featuresInQ8_leadingZeros_T_12063[25] ? 6'h19 :
    _featuresInQ8_leadingZeros_T_12134; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12136 = _featuresInQ8_leadingZeros_T_12063[24] ? 6'h18 :
    _featuresInQ8_leadingZeros_T_12135; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12137 = _featuresInQ8_leadingZeros_T_12063[23] ? 6'h17 :
    _featuresInQ8_leadingZeros_T_12136; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12138 = _featuresInQ8_leadingZeros_T_12063[22] ? 6'h16 :
    _featuresInQ8_leadingZeros_T_12137; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12139 = _featuresInQ8_leadingZeros_T_12063[21] ? 6'h15 :
    _featuresInQ8_leadingZeros_T_12138; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12140 = _featuresInQ8_leadingZeros_T_12063[20] ? 6'h14 :
    _featuresInQ8_leadingZeros_T_12139; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12141 = _featuresInQ8_leadingZeros_T_12063[19] ? 6'h13 :
    _featuresInQ8_leadingZeros_T_12140; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12142 = _featuresInQ8_leadingZeros_T_12063[18] ? 6'h12 :
    _featuresInQ8_leadingZeros_T_12141; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12143 = _featuresInQ8_leadingZeros_T_12063[17] ? 6'h11 :
    _featuresInQ8_leadingZeros_T_12142; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12144 = _featuresInQ8_leadingZeros_T_12063[16] ? 6'h10 :
    _featuresInQ8_leadingZeros_T_12143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12145 = _featuresInQ8_leadingZeros_T_12063[15] ? 6'hf :
    _featuresInQ8_leadingZeros_T_12144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12146 = _featuresInQ8_leadingZeros_T_12063[14] ? 6'he :
    _featuresInQ8_leadingZeros_T_12145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12147 = _featuresInQ8_leadingZeros_T_12063[13] ? 6'hd :
    _featuresInQ8_leadingZeros_T_12146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12148 = _featuresInQ8_leadingZeros_T_12063[12] ? 6'hc :
    _featuresInQ8_leadingZeros_T_12147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12149 = _featuresInQ8_leadingZeros_T_12063[11] ? 6'hb :
    _featuresInQ8_leadingZeros_T_12148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12150 = _featuresInQ8_leadingZeros_T_12063[10] ? 6'ha :
    _featuresInQ8_leadingZeros_T_12149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12151 = _featuresInQ8_leadingZeros_T_12063[9] ? 6'h9 :
    _featuresInQ8_leadingZeros_T_12150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12152 = _featuresInQ8_leadingZeros_T_12063[8] ? 6'h8 :
    _featuresInQ8_leadingZeros_T_12151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12153 = _featuresInQ8_leadingZeros_T_12063[7] ? 6'h7 :
    _featuresInQ8_leadingZeros_T_12152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12154 = _featuresInQ8_leadingZeros_T_12063[6] ? 6'h6 :
    _featuresInQ8_leadingZeros_T_12153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12155 = _featuresInQ8_leadingZeros_T_12063[5] ? 6'h5 :
    _featuresInQ8_leadingZeros_T_12154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12156 = _featuresInQ8_leadingZeros_T_12063[4] ? 6'h4 :
    _featuresInQ8_leadingZeros_T_12155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12157 = _featuresInQ8_leadingZeros_T_12063[3] ? 6'h3 :
    _featuresInQ8_leadingZeros_T_12156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12158 = _featuresInQ8_leadingZeros_T_12063[2] ? 6'h2 :
    _featuresInQ8_leadingZeros_T_12157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_leadingZeros_T_12159 = _featuresInQ8_leadingZeros_T_12063[1] ? 6'h1 :
    _featuresInQ8_leadingZeros_T_12158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] featuresInQ8_leadingZeros_63 = _featuresInQ8_leadingZeros_T_12063[0] ? 6'h0 :
    _featuresInQ8_leadingZeros_T_12159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _featuresInQ8_expRaw_T_127 = 6'h1f - featuresInQ8_leadingZeros_63; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] featuresInQ8_expRaw_63 = featuresInQ8_isZero_63 ? 6'h0 : _featuresInQ8_expRaw_T_127; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _featuresInQ8_shiftAmt_T_191 = featuresInQ8_expRaw_63 - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] featuresInQ8_shiftAmt_63 = featuresInQ8_expRaw_63 > 6'h3 ? _featuresInQ8_shiftAmt_T_191 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _featuresInQ8_mantissaRaw_T_63 = featuresInQ8_absClipped_63 >> featuresInQ8_shiftAmt_63; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] featuresInQ8_mantissaRaw_63 = _featuresInQ8_mantissaRaw_T_63[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] featuresInQ8_mantissa_63 = featuresInQ8_expRaw_63 >= 6'h3 ? featuresInQ8_mantissaRaw_63[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] featuresInQ8_expAdjusted_63 = featuresInQ8_expRaw_63 + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _featuresInQ8_exp_T_319 = featuresInQ8_expAdjusted_63 > 7'hf ? 4'hf : featuresInQ8_expAdjusted_63[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] featuresInQ8_exp_63 = featuresInQ8_isZero_63 ? 4'h0 : _featuresInQ8_exp_T_319; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] featuresInQ8_fp8_63 = {featuresInQ8_clippedX_63[31],featuresInQ8_exp_63,featuresInQ8_mantissa_63}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [7:0] featuresInQ8_63 = featuresInQ8_isZero_63 ? 8'h0 : featuresInQ8_fp8_63; // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
  reg [7:0] weightQ8_63_0; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_1; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_2; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_3; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_4; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_5; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_6; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_7; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_8; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_9; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_10; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_11; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_12; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_13; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_14; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_15; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_16; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_17; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_18; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_19; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_20; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_21; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_22; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_23; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_24; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_25; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_26; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_27; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_28; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_29; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_30; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  reg [7:0] weightQ8_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 115:23]
  wire [31:0] _weightQ8_63_0_T = {24'h0,linear_weight_63_0}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_0_sign = _weightQ8_63_0_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_0_absX_T = ~_weightQ8_63_0_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_0_absX_T_2 = _weightQ8_63_0_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_0_absX = weightQ8_63_0_sign ? _weightQ8_63_0_absX_T_2 : _weightQ8_63_0_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_0_shiftedX_T_1 = _GEN_14432 - weightQ8_63_0_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_0_shiftedX_T_3 = weightQ8_63_0_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_0_shiftedX = weightQ8_63_0_sign ? _weightQ8_63_0_shiftedX_T_1 : _weightQ8_63_0_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_0_scaledX_T_1 = weightQ8_63_0_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_0_scaledX = _weightQ8_63_0_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_0_clippedX_T_2 = weightQ8_63_0_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_0_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_0_clippedX = weightQ8_63_0_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_0_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_0_absClipped_T_1 = ~weightQ8_63_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_0_absClipped_T_3 = _weightQ8_63_0_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_0_absClipped = weightQ8_63_0_clippedX[31] ? _weightQ8_63_0_absClipped_T_3 :
    weightQ8_63_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_0_isZero = weightQ8_63_0_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37314 = {{16'd0}, weightQ8_63_0_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_4 = _GEN_37314 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_6 = {weightQ8_63_0_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_8 = _weightQ8_63_0_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_9 = _weightQ8_63_0_leadingZeros_T_4 | _weightQ8_63_0_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37315 = {{8'd0}, _weightQ8_63_0_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_14 = _GEN_37315 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_16 = {_weightQ8_63_0_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_18 = _weightQ8_63_0_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_19 = _weightQ8_63_0_leadingZeros_T_14 | _weightQ8_63_0_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37316 = {{4'd0}, _weightQ8_63_0_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_24 = _GEN_37316 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_26 = {_weightQ8_63_0_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_28 = _weightQ8_63_0_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_29 = _weightQ8_63_0_leadingZeros_T_24 | _weightQ8_63_0_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37317 = {{2'd0}, _weightQ8_63_0_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_34 = _GEN_37317 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_36 = {_weightQ8_63_0_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_38 = _weightQ8_63_0_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_39 = _weightQ8_63_0_leadingZeros_T_34 | _weightQ8_63_0_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37318 = {{1'd0}, _weightQ8_63_0_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_44 = _GEN_37318 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_46 = {_weightQ8_63_0_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_48 = _weightQ8_63_0_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_0_leadingZeros_T_49 = _weightQ8_63_0_leadingZeros_T_44 | _weightQ8_63_0_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37319 = {{8'd0}, weightQ8_63_0_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_55 = _GEN_37319 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_57 = {weightQ8_63_0_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_59 = _weightQ8_63_0_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_60 = _weightQ8_63_0_leadingZeros_T_55 | _weightQ8_63_0_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37320 = {{4'd0}, _weightQ8_63_0_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_65 = _GEN_37320 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_67 = {_weightQ8_63_0_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_69 = _weightQ8_63_0_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_70 = _weightQ8_63_0_leadingZeros_T_65 | _weightQ8_63_0_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37321 = {{2'd0}, _weightQ8_63_0_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_75 = _GEN_37321 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_77 = {_weightQ8_63_0_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_79 = _weightQ8_63_0_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_80 = _weightQ8_63_0_leadingZeros_T_75 | _weightQ8_63_0_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37322 = {{1'd0}, _weightQ8_63_0_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_85 = _GEN_37322 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_87 = {_weightQ8_63_0_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_89 = _weightQ8_63_0_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_0_leadingZeros_T_90 = _weightQ8_63_0_leadingZeros_T_85 | _weightQ8_63_0_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_0_leadingZeros_T_93 = {_weightQ8_63_0_leadingZeros_T_49,_weightQ8_63_0_leadingZeros_T_90,
    weightQ8_63_0_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_143 = _weightQ8_63_0_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_144 = _weightQ8_63_0_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_0_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_145 = _weightQ8_63_0_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_0_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_146 = _weightQ8_63_0_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_0_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_147 = _weightQ8_63_0_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_0_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_148 = _weightQ8_63_0_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_0_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_149 = _weightQ8_63_0_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_0_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_150 = _weightQ8_63_0_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_0_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_151 = _weightQ8_63_0_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_0_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_152 = _weightQ8_63_0_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_0_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_153 = _weightQ8_63_0_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_0_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_154 = _weightQ8_63_0_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_0_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_155 = _weightQ8_63_0_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_0_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_156 = _weightQ8_63_0_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_0_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_157 = _weightQ8_63_0_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_0_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_158 = _weightQ8_63_0_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_0_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_159 = _weightQ8_63_0_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_0_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_160 = _weightQ8_63_0_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_0_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_161 = _weightQ8_63_0_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_0_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_162 = _weightQ8_63_0_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_0_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_163 = _weightQ8_63_0_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_0_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_164 = _weightQ8_63_0_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_0_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_165 = _weightQ8_63_0_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_0_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_166 = _weightQ8_63_0_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_0_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_167 = _weightQ8_63_0_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_0_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_168 = _weightQ8_63_0_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_0_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_169 = _weightQ8_63_0_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_0_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_170 = _weightQ8_63_0_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_0_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_171 = _weightQ8_63_0_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_0_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_172 = _weightQ8_63_0_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_0_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_173 = _weightQ8_63_0_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_0_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_174 = _weightQ8_63_0_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_0_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_175 = _weightQ8_63_0_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_0_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_176 = _weightQ8_63_0_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_0_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_177 = _weightQ8_63_0_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_0_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_178 = _weightQ8_63_0_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_0_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_179 = _weightQ8_63_0_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_0_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_180 = _weightQ8_63_0_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_0_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_181 = _weightQ8_63_0_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_0_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_182 = _weightQ8_63_0_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_0_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_183 = _weightQ8_63_0_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_0_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_184 = _weightQ8_63_0_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_0_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_185 = _weightQ8_63_0_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_0_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_186 = _weightQ8_63_0_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_0_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_187 = _weightQ8_63_0_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_0_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_188 = _weightQ8_63_0_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_0_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_leadingZeros_T_189 = _weightQ8_63_0_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_0_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_0_leadingZeros = _weightQ8_63_0_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_0_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_0_expRaw_T_1 = 6'h1f - weightQ8_63_0_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_0_expRaw = weightQ8_63_0_isZero ? 6'h0 : _weightQ8_63_0_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_0_shiftAmt_T_2 = weightQ8_63_0_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_0_shiftAmt = weightQ8_63_0_expRaw > 6'h3 ? _weightQ8_63_0_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_0_mantissaRaw_T = weightQ8_63_0_absClipped >> weightQ8_63_0_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_0_mantissaRaw = _weightQ8_63_0_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_0_mantissa = weightQ8_63_0_expRaw >= 6'h3 ? weightQ8_63_0_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_0_expAdjusted = weightQ8_63_0_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_0_exp_T_4 = weightQ8_63_0_expAdjusted > 7'hf ? 4'hf : weightQ8_63_0_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_0_exp = weightQ8_63_0_isZero ? 4'h0 : _weightQ8_63_0_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_0_fp8 = {weightQ8_63_0_clippedX[31],weightQ8_63_0_exp,weightQ8_63_0_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_1_T = {24'h0,linear_weight_63_1}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_1_sign = _weightQ8_63_1_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_1_absX_T = ~_weightQ8_63_1_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_1_absX_T_2 = _weightQ8_63_1_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_1_absX = weightQ8_63_1_sign ? _weightQ8_63_1_absX_T_2 : _weightQ8_63_1_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_1_shiftedX_T_1 = _GEN_14432 - weightQ8_63_1_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_1_shiftedX_T_3 = weightQ8_63_1_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_1_shiftedX = weightQ8_63_1_sign ? _weightQ8_63_1_shiftedX_T_1 : _weightQ8_63_1_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_1_scaledX_T_1 = weightQ8_63_1_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_1_scaledX = _weightQ8_63_1_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_1_clippedX_T_2 = weightQ8_63_1_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_1_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_1_clippedX = weightQ8_63_1_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_1_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_1_absClipped_T_1 = ~weightQ8_63_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_1_absClipped_T_3 = _weightQ8_63_1_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_1_absClipped = weightQ8_63_1_clippedX[31] ? _weightQ8_63_1_absClipped_T_3 :
    weightQ8_63_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_1_isZero = weightQ8_63_1_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37325 = {{16'd0}, weightQ8_63_1_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_4 = _GEN_37325 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_6 = {weightQ8_63_1_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_8 = _weightQ8_63_1_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_9 = _weightQ8_63_1_leadingZeros_T_4 | _weightQ8_63_1_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37326 = {{8'd0}, _weightQ8_63_1_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_14 = _GEN_37326 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_16 = {_weightQ8_63_1_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_18 = _weightQ8_63_1_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_19 = _weightQ8_63_1_leadingZeros_T_14 | _weightQ8_63_1_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37327 = {{4'd0}, _weightQ8_63_1_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_24 = _GEN_37327 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_26 = {_weightQ8_63_1_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_28 = _weightQ8_63_1_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_29 = _weightQ8_63_1_leadingZeros_T_24 | _weightQ8_63_1_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37328 = {{2'd0}, _weightQ8_63_1_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_34 = _GEN_37328 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_36 = {_weightQ8_63_1_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_38 = _weightQ8_63_1_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_39 = _weightQ8_63_1_leadingZeros_T_34 | _weightQ8_63_1_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37329 = {{1'd0}, _weightQ8_63_1_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_44 = _GEN_37329 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_46 = {_weightQ8_63_1_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_48 = _weightQ8_63_1_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_1_leadingZeros_T_49 = _weightQ8_63_1_leadingZeros_T_44 | _weightQ8_63_1_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37330 = {{8'd0}, weightQ8_63_1_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_55 = _GEN_37330 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_57 = {weightQ8_63_1_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_59 = _weightQ8_63_1_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_60 = _weightQ8_63_1_leadingZeros_T_55 | _weightQ8_63_1_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37331 = {{4'd0}, _weightQ8_63_1_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_65 = _GEN_37331 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_67 = {_weightQ8_63_1_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_69 = _weightQ8_63_1_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_70 = _weightQ8_63_1_leadingZeros_T_65 | _weightQ8_63_1_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37332 = {{2'd0}, _weightQ8_63_1_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_75 = _GEN_37332 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_77 = {_weightQ8_63_1_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_79 = _weightQ8_63_1_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_80 = _weightQ8_63_1_leadingZeros_T_75 | _weightQ8_63_1_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37333 = {{1'd0}, _weightQ8_63_1_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_85 = _GEN_37333 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_87 = {_weightQ8_63_1_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_89 = _weightQ8_63_1_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_1_leadingZeros_T_90 = _weightQ8_63_1_leadingZeros_T_85 | _weightQ8_63_1_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_1_leadingZeros_T_93 = {_weightQ8_63_1_leadingZeros_T_49,_weightQ8_63_1_leadingZeros_T_90,
    weightQ8_63_1_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_143 = _weightQ8_63_1_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_144 = _weightQ8_63_1_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_1_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_145 = _weightQ8_63_1_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_1_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_146 = _weightQ8_63_1_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_1_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_147 = _weightQ8_63_1_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_1_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_148 = _weightQ8_63_1_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_1_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_149 = _weightQ8_63_1_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_1_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_150 = _weightQ8_63_1_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_1_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_151 = _weightQ8_63_1_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_1_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_152 = _weightQ8_63_1_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_1_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_153 = _weightQ8_63_1_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_1_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_154 = _weightQ8_63_1_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_1_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_155 = _weightQ8_63_1_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_1_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_156 = _weightQ8_63_1_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_1_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_157 = _weightQ8_63_1_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_1_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_158 = _weightQ8_63_1_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_1_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_159 = _weightQ8_63_1_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_1_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_160 = _weightQ8_63_1_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_1_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_161 = _weightQ8_63_1_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_1_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_162 = _weightQ8_63_1_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_1_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_163 = _weightQ8_63_1_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_1_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_164 = _weightQ8_63_1_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_1_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_165 = _weightQ8_63_1_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_1_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_166 = _weightQ8_63_1_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_1_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_167 = _weightQ8_63_1_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_1_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_168 = _weightQ8_63_1_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_1_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_169 = _weightQ8_63_1_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_1_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_170 = _weightQ8_63_1_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_1_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_171 = _weightQ8_63_1_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_1_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_172 = _weightQ8_63_1_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_1_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_173 = _weightQ8_63_1_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_1_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_174 = _weightQ8_63_1_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_1_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_175 = _weightQ8_63_1_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_1_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_176 = _weightQ8_63_1_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_1_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_177 = _weightQ8_63_1_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_1_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_178 = _weightQ8_63_1_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_1_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_179 = _weightQ8_63_1_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_1_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_180 = _weightQ8_63_1_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_1_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_181 = _weightQ8_63_1_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_1_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_182 = _weightQ8_63_1_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_1_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_183 = _weightQ8_63_1_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_1_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_184 = _weightQ8_63_1_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_1_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_185 = _weightQ8_63_1_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_1_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_186 = _weightQ8_63_1_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_1_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_187 = _weightQ8_63_1_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_1_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_188 = _weightQ8_63_1_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_1_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_leadingZeros_T_189 = _weightQ8_63_1_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_1_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_1_leadingZeros = _weightQ8_63_1_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_1_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_1_expRaw_T_1 = 6'h1f - weightQ8_63_1_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_1_expRaw = weightQ8_63_1_isZero ? 6'h0 : _weightQ8_63_1_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_1_shiftAmt_T_2 = weightQ8_63_1_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_1_shiftAmt = weightQ8_63_1_expRaw > 6'h3 ? _weightQ8_63_1_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_1_mantissaRaw_T = weightQ8_63_1_absClipped >> weightQ8_63_1_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_1_mantissaRaw = _weightQ8_63_1_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_1_mantissa = weightQ8_63_1_expRaw >= 6'h3 ? weightQ8_63_1_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_1_expAdjusted = weightQ8_63_1_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_1_exp_T_4 = weightQ8_63_1_expAdjusted > 7'hf ? 4'hf : weightQ8_63_1_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_1_exp = weightQ8_63_1_isZero ? 4'h0 : _weightQ8_63_1_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_1_fp8 = {weightQ8_63_1_clippedX[31],weightQ8_63_1_exp,weightQ8_63_1_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_2_T = {24'h0,linear_weight_63_2}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_2_sign = _weightQ8_63_2_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_2_absX_T = ~_weightQ8_63_2_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_2_absX_T_2 = _weightQ8_63_2_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_2_absX = weightQ8_63_2_sign ? _weightQ8_63_2_absX_T_2 : _weightQ8_63_2_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_2_shiftedX_T_1 = _GEN_14432 - weightQ8_63_2_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_2_shiftedX_T_3 = weightQ8_63_2_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_2_shiftedX = weightQ8_63_2_sign ? _weightQ8_63_2_shiftedX_T_1 : _weightQ8_63_2_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_2_scaledX_T_1 = weightQ8_63_2_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_2_scaledX = _weightQ8_63_2_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_2_clippedX_T_2 = weightQ8_63_2_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_2_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_2_clippedX = weightQ8_63_2_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_2_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_2_absClipped_T_1 = ~weightQ8_63_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_2_absClipped_T_3 = _weightQ8_63_2_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_2_absClipped = weightQ8_63_2_clippedX[31] ? _weightQ8_63_2_absClipped_T_3 :
    weightQ8_63_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_2_isZero = weightQ8_63_2_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37336 = {{16'd0}, weightQ8_63_2_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_4 = _GEN_37336 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_6 = {weightQ8_63_2_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_8 = _weightQ8_63_2_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_9 = _weightQ8_63_2_leadingZeros_T_4 | _weightQ8_63_2_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37337 = {{8'd0}, _weightQ8_63_2_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_14 = _GEN_37337 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_16 = {_weightQ8_63_2_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_18 = _weightQ8_63_2_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_19 = _weightQ8_63_2_leadingZeros_T_14 | _weightQ8_63_2_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37338 = {{4'd0}, _weightQ8_63_2_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_24 = _GEN_37338 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_26 = {_weightQ8_63_2_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_28 = _weightQ8_63_2_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_29 = _weightQ8_63_2_leadingZeros_T_24 | _weightQ8_63_2_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37339 = {{2'd0}, _weightQ8_63_2_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_34 = _GEN_37339 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_36 = {_weightQ8_63_2_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_38 = _weightQ8_63_2_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_39 = _weightQ8_63_2_leadingZeros_T_34 | _weightQ8_63_2_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37340 = {{1'd0}, _weightQ8_63_2_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_44 = _GEN_37340 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_46 = {_weightQ8_63_2_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_48 = _weightQ8_63_2_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_2_leadingZeros_T_49 = _weightQ8_63_2_leadingZeros_T_44 | _weightQ8_63_2_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37341 = {{8'd0}, weightQ8_63_2_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_55 = _GEN_37341 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_57 = {weightQ8_63_2_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_59 = _weightQ8_63_2_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_60 = _weightQ8_63_2_leadingZeros_T_55 | _weightQ8_63_2_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37342 = {{4'd0}, _weightQ8_63_2_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_65 = _GEN_37342 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_67 = {_weightQ8_63_2_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_69 = _weightQ8_63_2_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_70 = _weightQ8_63_2_leadingZeros_T_65 | _weightQ8_63_2_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37343 = {{2'd0}, _weightQ8_63_2_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_75 = _GEN_37343 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_77 = {_weightQ8_63_2_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_79 = _weightQ8_63_2_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_80 = _weightQ8_63_2_leadingZeros_T_75 | _weightQ8_63_2_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37344 = {{1'd0}, _weightQ8_63_2_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_85 = _GEN_37344 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_87 = {_weightQ8_63_2_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_89 = _weightQ8_63_2_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_2_leadingZeros_T_90 = _weightQ8_63_2_leadingZeros_T_85 | _weightQ8_63_2_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_2_leadingZeros_T_93 = {_weightQ8_63_2_leadingZeros_T_49,_weightQ8_63_2_leadingZeros_T_90,
    weightQ8_63_2_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_143 = _weightQ8_63_2_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_144 = _weightQ8_63_2_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_2_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_145 = _weightQ8_63_2_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_2_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_146 = _weightQ8_63_2_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_2_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_147 = _weightQ8_63_2_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_2_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_148 = _weightQ8_63_2_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_2_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_149 = _weightQ8_63_2_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_2_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_150 = _weightQ8_63_2_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_2_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_151 = _weightQ8_63_2_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_2_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_152 = _weightQ8_63_2_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_2_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_153 = _weightQ8_63_2_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_2_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_154 = _weightQ8_63_2_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_2_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_155 = _weightQ8_63_2_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_2_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_156 = _weightQ8_63_2_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_2_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_157 = _weightQ8_63_2_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_2_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_158 = _weightQ8_63_2_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_2_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_159 = _weightQ8_63_2_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_2_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_160 = _weightQ8_63_2_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_2_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_161 = _weightQ8_63_2_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_2_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_162 = _weightQ8_63_2_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_2_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_163 = _weightQ8_63_2_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_2_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_164 = _weightQ8_63_2_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_2_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_165 = _weightQ8_63_2_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_2_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_166 = _weightQ8_63_2_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_2_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_167 = _weightQ8_63_2_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_2_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_168 = _weightQ8_63_2_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_2_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_169 = _weightQ8_63_2_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_2_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_170 = _weightQ8_63_2_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_2_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_171 = _weightQ8_63_2_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_2_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_172 = _weightQ8_63_2_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_2_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_173 = _weightQ8_63_2_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_2_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_174 = _weightQ8_63_2_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_2_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_175 = _weightQ8_63_2_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_2_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_176 = _weightQ8_63_2_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_2_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_177 = _weightQ8_63_2_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_2_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_178 = _weightQ8_63_2_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_2_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_179 = _weightQ8_63_2_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_2_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_180 = _weightQ8_63_2_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_2_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_181 = _weightQ8_63_2_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_2_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_182 = _weightQ8_63_2_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_2_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_183 = _weightQ8_63_2_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_2_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_184 = _weightQ8_63_2_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_2_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_185 = _weightQ8_63_2_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_2_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_186 = _weightQ8_63_2_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_2_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_187 = _weightQ8_63_2_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_2_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_188 = _weightQ8_63_2_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_2_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_leadingZeros_T_189 = _weightQ8_63_2_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_2_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_2_leadingZeros = _weightQ8_63_2_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_2_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_2_expRaw_T_1 = 6'h1f - weightQ8_63_2_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_2_expRaw = weightQ8_63_2_isZero ? 6'h0 : _weightQ8_63_2_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_2_shiftAmt_T_2 = weightQ8_63_2_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_2_shiftAmt = weightQ8_63_2_expRaw > 6'h3 ? _weightQ8_63_2_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_2_mantissaRaw_T = weightQ8_63_2_absClipped >> weightQ8_63_2_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_2_mantissaRaw = _weightQ8_63_2_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_2_mantissa = weightQ8_63_2_expRaw >= 6'h3 ? weightQ8_63_2_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_2_expAdjusted = weightQ8_63_2_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_2_exp_T_4 = weightQ8_63_2_expAdjusted > 7'hf ? 4'hf : weightQ8_63_2_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_2_exp = weightQ8_63_2_isZero ? 4'h0 : _weightQ8_63_2_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_2_fp8 = {weightQ8_63_2_clippedX[31],weightQ8_63_2_exp,weightQ8_63_2_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_3_T = {24'h0,linear_weight_63_3}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_3_sign = _weightQ8_63_3_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_3_absX_T = ~_weightQ8_63_3_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_3_absX_T_2 = _weightQ8_63_3_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_3_absX = weightQ8_63_3_sign ? _weightQ8_63_3_absX_T_2 : _weightQ8_63_3_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_3_shiftedX_T_1 = _GEN_14432 - weightQ8_63_3_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_3_shiftedX_T_3 = weightQ8_63_3_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_3_shiftedX = weightQ8_63_3_sign ? _weightQ8_63_3_shiftedX_T_1 : _weightQ8_63_3_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_3_scaledX_T_1 = weightQ8_63_3_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_3_scaledX = _weightQ8_63_3_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_3_clippedX_T_2 = weightQ8_63_3_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_3_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_3_clippedX = weightQ8_63_3_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_3_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_3_absClipped_T_1 = ~weightQ8_63_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_3_absClipped_T_3 = _weightQ8_63_3_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_3_absClipped = weightQ8_63_3_clippedX[31] ? _weightQ8_63_3_absClipped_T_3 :
    weightQ8_63_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_3_isZero = weightQ8_63_3_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37347 = {{16'd0}, weightQ8_63_3_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_4 = _GEN_37347 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_6 = {weightQ8_63_3_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_8 = _weightQ8_63_3_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_9 = _weightQ8_63_3_leadingZeros_T_4 | _weightQ8_63_3_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37348 = {{8'd0}, _weightQ8_63_3_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_14 = _GEN_37348 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_16 = {_weightQ8_63_3_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_18 = _weightQ8_63_3_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_19 = _weightQ8_63_3_leadingZeros_T_14 | _weightQ8_63_3_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37349 = {{4'd0}, _weightQ8_63_3_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_24 = _GEN_37349 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_26 = {_weightQ8_63_3_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_28 = _weightQ8_63_3_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_29 = _weightQ8_63_3_leadingZeros_T_24 | _weightQ8_63_3_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37350 = {{2'd0}, _weightQ8_63_3_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_34 = _GEN_37350 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_36 = {_weightQ8_63_3_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_38 = _weightQ8_63_3_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_39 = _weightQ8_63_3_leadingZeros_T_34 | _weightQ8_63_3_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37351 = {{1'd0}, _weightQ8_63_3_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_44 = _GEN_37351 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_46 = {_weightQ8_63_3_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_48 = _weightQ8_63_3_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_3_leadingZeros_T_49 = _weightQ8_63_3_leadingZeros_T_44 | _weightQ8_63_3_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37352 = {{8'd0}, weightQ8_63_3_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_55 = _GEN_37352 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_57 = {weightQ8_63_3_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_59 = _weightQ8_63_3_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_60 = _weightQ8_63_3_leadingZeros_T_55 | _weightQ8_63_3_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37353 = {{4'd0}, _weightQ8_63_3_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_65 = _GEN_37353 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_67 = {_weightQ8_63_3_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_69 = _weightQ8_63_3_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_70 = _weightQ8_63_3_leadingZeros_T_65 | _weightQ8_63_3_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37354 = {{2'd0}, _weightQ8_63_3_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_75 = _GEN_37354 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_77 = {_weightQ8_63_3_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_79 = _weightQ8_63_3_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_80 = _weightQ8_63_3_leadingZeros_T_75 | _weightQ8_63_3_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37355 = {{1'd0}, _weightQ8_63_3_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_85 = _GEN_37355 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_87 = {_weightQ8_63_3_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_89 = _weightQ8_63_3_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_3_leadingZeros_T_90 = _weightQ8_63_3_leadingZeros_T_85 | _weightQ8_63_3_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_3_leadingZeros_T_93 = {_weightQ8_63_3_leadingZeros_T_49,_weightQ8_63_3_leadingZeros_T_90,
    weightQ8_63_3_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_143 = _weightQ8_63_3_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_144 = _weightQ8_63_3_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_3_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_145 = _weightQ8_63_3_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_3_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_146 = _weightQ8_63_3_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_3_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_147 = _weightQ8_63_3_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_3_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_148 = _weightQ8_63_3_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_3_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_149 = _weightQ8_63_3_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_3_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_150 = _weightQ8_63_3_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_3_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_151 = _weightQ8_63_3_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_3_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_152 = _weightQ8_63_3_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_3_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_153 = _weightQ8_63_3_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_3_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_154 = _weightQ8_63_3_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_3_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_155 = _weightQ8_63_3_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_3_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_156 = _weightQ8_63_3_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_3_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_157 = _weightQ8_63_3_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_3_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_158 = _weightQ8_63_3_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_3_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_159 = _weightQ8_63_3_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_3_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_160 = _weightQ8_63_3_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_3_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_161 = _weightQ8_63_3_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_3_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_162 = _weightQ8_63_3_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_3_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_163 = _weightQ8_63_3_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_3_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_164 = _weightQ8_63_3_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_3_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_165 = _weightQ8_63_3_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_3_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_166 = _weightQ8_63_3_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_3_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_167 = _weightQ8_63_3_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_3_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_168 = _weightQ8_63_3_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_3_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_169 = _weightQ8_63_3_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_3_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_170 = _weightQ8_63_3_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_3_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_171 = _weightQ8_63_3_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_3_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_172 = _weightQ8_63_3_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_3_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_173 = _weightQ8_63_3_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_3_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_174 = _weightQ8_63_3_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_3_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_175 = _weightQ8_63_3_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_3_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_176 = _weightQ8_63_3_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_3_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_177 = _weightQ8_63_3_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_3_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_178 = _weightQ8_63_3_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_3_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_179 = _weightQ8_63_3_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_3_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_180 = _weightQ8_63_3_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_3_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_181 = _weightQ8_63_3_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_3_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_182 = _weightQ8_63_3_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_3_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_183 = _weightQ8_63_3_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_3_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_184 = _weightQ8_63_3_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_3_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_185 = _weightQ8_63_3_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_3_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_186 = _weightQ8_63_3_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_3_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_187 = _weightQ8_63_3_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_3_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_188 = _weightQ8_63_3_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_3_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_leadingZeros_T_189 = _weightQ8_63_3_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_3_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_3_leadingZeros = _weightQ8_63_3_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_3_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_3_expRaw_T_1 = 6'h1f - weightQ8_63_3_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_3_expRaw = weightQ8_63_3_isZero ? 6'h0 : _weightQ8_63_3_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_3_shiftAmt_T_2 = weightQ8_63_3_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_3_shiftAmt = weightQ8_63_3_expRaw > 6'h3 ? _weightQ8_63_3_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_3_mantissaRaw_T = weightQ8_63_3_absClipped >> weightQ8_63_3_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_3_mantissaRaw = _weightQ8_63_3_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_3_mantissa = weightQ8_63_3_expRaw >= 6'h3 ? weightQ8_63_3_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_3_expAdjusted = weightQ8_63_3_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_3_exp_T_4 = weightQ8_63_3_expAdjusted > 7'hf ? 4'hf : weightQ8_63_3_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_3_exp = weightQ8_63_3_isZero ? 4'h0 : _weightQ8_63_3_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_3_fp8 = {weightQ8_63_3_clippedX[31],weightQ8_63_3_exp,weightQ8_63_3_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_4_T = {24'h0,linear_weight_63_4}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_4_sign = _weightQ8_63_4_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_4_absX_T = ~_weightQ8_63_4_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_4_absX_T_2 = _weightQ8_63_4_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_4_absX = weightQ8_63_4_sign ? _weightQ8_63_4_absX_T_2 : _weightQ8_63_4_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_4_shiftedX_T_1 = _GEN_14432 - weightQ8_63_4_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_4_shiftedX_T_3 = weightQ8_63_4_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_4_shiftedX = weightQ8_63_4_sign ? _weightQ8_63_4_shiftedX_T_1 : _weightQ8_63_4_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_4_scaledX_T_1 = weightQ8_63_4_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_4_scaledX = _weightQ8_63_4_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_4_clippedX_T_2 = weightQ8_63_4_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_4_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_4_clippedX = weightQ8_63_4_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_4_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_4_absClipped_T_1 = ~weightQ8_63_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_4_absClipped_T_3 = _weightQ8_63_4_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_4_absClipped = weightQ8_63_4_clippedX[31] ? _weightQ8_63_4_absClipped_T_3 :
    weightQ8_63_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_4_isZero = weightQ8_63_4_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37358 = {{16'd0}, weightQ8_63_4_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_4 = _GEN_37358 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_6 = {weightQ8_63_4_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_8 = _weightQ8_63_4_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_9 = _weightQ8_63_4_leadingZeros_T_4 | _weightQ8_63_4_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37359 = {{8'd0}, _weightQ8_63_4_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_14 = _GEN_37359 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_16 = {_weightQ8_63_4_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_18 = _weightQ8_63_4_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_19 = _weightQ8_63_4_leadingZeros_T_14 | _weightQ8_63_4_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37360 = {{4'd0}, _weightQ8_63_4_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_24 = _GEN_37360 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_26 = {_weightQ8_63_4_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_28 = _weightQ8_63_4_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_29 = _weightQ8_63_4_leadingZeros_T_24 | _weightQ8_63_4_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37361 = {{2'd0}, _weightQ8_63_4_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_34 = _GEN_37361 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_36 = {_weightQ8_63_4_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_38 = _weightQ8_63_4_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_39 = _weightQ8_63_4_leadingZeros_T_34 | _weightQ8_63_4_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37362 = {{1'd0}, _weightQ8_63_4_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_44 = _GEN_37362 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_46 = {_weightQ8_63_4_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_48 = _weightQ8_63_4_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_4_leadingZeros_T_49 = _weightQ8_63_4_leadingZeros_T_44 | _weightQ8_63_4_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37363 = {{8'd0}, weightQ8_63_4_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_55 = _GEN_37363 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_57 = {weightQ8_63_4_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_59 = _weightQ8_63_4_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_60 = _weightQ8_63_4_leadingZeros_T_55 | _weightQ8_63_4_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37364 = {{4'd0}, _weightQ8_63_4_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_65 = _GEN_37364 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_67 = {_weightQ8_63_4_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_69 = _weightQ8_63_4_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_70 = _weightQ8_63_4_leadingZeros_T_65 | _weightQ8_63_4_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37365 = {{2'd0}, _weightQ8_63_4_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_75 = _GEN_37365 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_77 = {_weightQ8_63_4_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_79 = _weightQ8_63_4_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_80 = _weightQ8_63_4_leadingZeros_T_75 | _weightQ8_63_4_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37366 = {{1'd0}, _weightQ8_63_4_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_85 = _GEN_37366 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_87 = {_weightQ8_63_4_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_89 = _weightQ8_63_4_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_4_leadingZeros_T_90 = _weightQ8_63_4_leadingZeros_T_85 | _weightQ8_63_4_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_4_leadingZeros_T_93 = {_weightQ8_63_4_leadingZeros_T_49,_weightQ8_63_4_leadingZeros_T_90,
    weightQ8_63_4_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_143 = _weightQ8_63_4_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_144 = _weightQ8_63_4_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_4_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_145 = _weightQ8_63_4_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_4_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_146 = _weightQ8_63_4_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_4_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_147 = _weightQ8_63_4_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_4_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_148 = _weightQ8_63_4_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_4_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_149 = _weightQ8_63_4_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_4_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_150 = _weightQ8_63_4_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_4_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_151 = _weightQ8_63_4_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_4_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_152 = _weightQ8_63_4_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_4_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_153 = _weightQ8_63_4_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_4_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_154 = _weightQ8_63_4_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_4_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_155 = _weightQ8_63_4_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_4_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_156 = _weightQ8_63_4_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_4_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_157 = _weightQ8_63_4_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_4_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_158 = _weightQ8_63_4_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_4_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_159 = _weightQ8_63_4_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_4_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_160 = _weightQ8_63_4_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_4_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_161 = _weightQ8_63_4_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_4_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_162 = _weightQ8_63_4_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_4_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_163 = _weightQ8_63_4_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_4_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_164 = _weightQ8_63_4_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_4_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_165 = _weightQ8_63_4_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_4_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_166 = _weightQ8_63_4_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_4_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_167 = _weightQ8_63_4_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_4_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_168 = _weightQ8_63_4_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_4_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_169 = _weightQ8_63_4_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_4_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_170 = _weightQ8_63_4_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_4_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_171 = _weightQ8_63_4_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_4_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_172 = _weightQ8_63_4_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_4_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_173 = _weightQ8_63_4_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_4_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_174 = _weightQ8_63_4_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_4_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_175 = _weightQ8_63_4_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_4_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_176 = _weightQ8_63_4_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_4_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_177 = _weightQ8_63_4_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_4_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_178 = _weightQ8_63_4_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_4_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_179 = _weightQ8_63_4_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_4_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_180 = _weightQ8_63_4_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_4_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_181 = _weightQ8_63_4_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_4_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_182 = _weightQ8_63_4_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_4_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_183 = _weightQ8_63_4_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_4_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_184 = _weightQ8_63_4_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_4_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_185 = _weightQ8_63_4_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_4_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_186 = _weightQ8_63_4_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_4_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_187 = _weightQ8_63_4_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_4_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_188 = _weightQ8_63_4_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_4_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_leadingZeros_T_189 = _weightQ8_63_4_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_4_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_4_leadingZeros = _weightQ8_63_4_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_4_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_4_expRaw_T_1 = 6'h1f - weightQ8_63_4_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_4_expRaw = weightQ8_63_4_isZero ? 6'h0 : _weightQ8_63_4_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_4_shiftAmt_T_2 = weightQ8_63_4_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_4_shiftAmt = weightQ8_63_4_expRaw > 6'h3 ? _weightQ8_63_4_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_4_mantissaRaw_T = weightQ8_63_4_absClipped >> weightQ8_63_4_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_4_mantissaRaw = _weightQ8_63_4_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_4_mantissa = weightQ8_63_4_expRaw >= 6'h3 ? weightQ8_63_4_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_4_expAdjusted = weightQ8_63_4_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_4_exp_T_4 = weightQ8_63_4_expAdjusted > 7'hf ? 4'hf : weightQ8_63_4_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_4_exp = weightQ8_63_4_isZero ? 4'h0 : _weightQ8_63_4_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_4_fp8 = {weightQ8_63_4_clippedX[31],weightQ8_63_4_exp,weightQ8_63_4_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_5_T = {24'h0,linear_weight_63_5}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_5_sign = _weightQ8_63_5_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_5_absX_T = ~_weightQ8_63_5_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_5_absX_T_2 = _weightQ8_63_5_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_5_absX = weightQ8_63_5_sign ? _weightQ8_63_5_absX_T_2 : _weightQ8_63_5_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_5_shiftedX_T_1 = _GEN_14432 - weightQ8_63_5_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_5_shiftedX_T_3 = weightQ8_63_5_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_5_shiftedX = weightQ8_63_5_sign ? _weightQ8_63_5_shiftedX_T_1 : _weightQ8_63_5_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_5_scaledX_T_1 = weightQ8_63_5_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_5_scaledX = _weightQ8_63_5_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_5_clippedX_T_2 = weightQ8_63_5_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_5_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_5_clippedX = weightQ8_63_5_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_5_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_5_absClipped_T_1 = ~weightQ8_63_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_5_absClipped_T_3 = _weightQ8_63_5_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_5_absClipped = weightQ8_63_5_clippedX[31] ? _weightQ8_63_5_absClipped_T_3 :
    weightQ8_63_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_5_isZero = weightQ8_63_5_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37369 = {{16'd0}, weightQ8_63_5_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_4 = _GEN_37369 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_6 = {weightQ8_63_5_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_8 = _weightQ8_63_5_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_9 = _weightQ8_63_5_leadingZeros_T_4 | _weightQ8_63_5_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37370 = {{8'd0}, _weightQ8_63_5_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_14 = _GEN_37370 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_16 = {_weightQ8_63_5_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_18 = _weightQ8_63_5_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_19 = _weightQ8_63_5_leadingZeros_T_14 | _weightQ8_63_5_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37371 = {{4'd0}, _weightQ8_63_5_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_24 = _GEN_37371 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_26 = {_weightQ8_63_5_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_28 = _weightQ8_63_5_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_29 = _weightQ8_63_5_leadingZeros_T_24 | _weightQ8_63_5_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37372 = {{2'd0}, _weightQ8_63_5_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_34 = _GEN_37372 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_36 = {_weightQ8_63_5_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_38 = _weightQ8_63_5_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_39 = _weightQ8_63_5_leadingZeros_T_34 | _weightQ8_63_5_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37373 = {{1'd0}, _weightQ8_63_5_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_44 = _GEN_37373 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_46 = {_weightQ8_63_5_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_48 = _weightQ8_63_5_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_5_leadingZeros_T_49 = _weightQ8_63_5_leadingZeros_T_44 | _weightQ8_63_5_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37374 = {{8'd0}, weightQ8_63_5_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_55 = _GEN_37374 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_57 = {weightQ8_63_5_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_59 = _weightQ8_63_5_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_60 = _weightQ8_63_5_leadingZeros_T_55 | _weightQ8_63_5_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37375 = {{4'd0}, _weightQ8_63_5_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_65 = _GEN_37375 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_67 = {_weightQ8_63_5_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_69 = _weightQ8_63_5_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_70 = _weightQ8_63_5_leadingZeros_T_65 | _weightQ8_63_5_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37376 = {{2'd0}, _weightQ8_63_5_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_75 = _GEN_37376 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_77 = {_weightQ8_63_5_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_79 = _weightQ8_63_5_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_80 = _weightQ8_63_5_leadingZeros_T_75 | _weightQ8_63_5_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37377 = {{1'd0}, _weightQ8_63_5_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_85 = _GEN_37377 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_87 = {_weightQ8_63_5_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_89 = _weightQ8_63_5_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_5_leadingZeros_T_90 = _weightQ8_63_5_leadingZeros_T_85 | _weightQ8_63_5_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_5_leadingZeros_T_93 = {_weightQ8_63_5_leadingZeros_T_49,_weightQ8_63_5_leadingZeros_T_90,
    weightQ8_63_5_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_143 = _weightQ8_63_5_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_144 = _weightQ8_63_5_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_5_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_145 = _weightQ8_63_5_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_5_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_146 = _weightQ8_63_5_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_5_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_147 = _weightQ8_63_5_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_5_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_148 = _weightQ8_63_5_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_5_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_149 = _weightQ8_63_5_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_5_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_150 = _weightQ8_63_5_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_5_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_151 = _weightQ8_63_5_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_5_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_152 = _weightQ8_63_5_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_5_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_153 = _weightQ8_63_5_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_5_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_154 = _weightQ8_63_5_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_5_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_155 = _weightQ8_63_5_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_5_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_156 = _weightQ8_63_5_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_5_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_157 = _weightQ8_63_5_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_5_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_158 = _weightQ8_63_5_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_5_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_159 = _weightQ8_63_5_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_5_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_160 = _weightQ8_63_5_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_5_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_161 = _weightQ8_63_5_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_5_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_162 = _weightQ8_63_5_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_5_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_163 = _weightQ8_63_5_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_5_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_164 = _weightQ8_63_5_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_5_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_165 = _weightQ8_63_5_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_5_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_166 = _weightQ8_63_5_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_5_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_167 = _weightQ8_63_5_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_5_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_168 = _weightQ8_63_5_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_5_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_169 = _weightQ8_63_5_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_5_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_170 = _weightQ8_63_5_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_5_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_171 = _weightQ8_63_5_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_5_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_172 = _weightQ8_63_5_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_5_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_173 = _weightQ8_63_5_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_5_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_174 = _weightQ8_63_5_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_5_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_175 = _weightQ8_63_5_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_5_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_176 = _weightQ8_63_5_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_5_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_177 = _weightQ8_63_5_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_5_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_178 = _weightQ8_63_5_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_5_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_179 = _weightQ8_63_5_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_5_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_180 = _weightQ8_63_5_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_5_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_181 = _weightQ8_63_5_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_5_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_182 = _weightQ8_63_5_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_5_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_183 = _weightQ8_63_5_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_5_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_184 = _weightQ8_63_5_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_5_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_185 = _weightQ8_63_5_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_5_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_186 = _weightQ8_63_5_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_5_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_187 = _weightQ8_63_5_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_5_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_188 = _weightQ8_63_5_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_5_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_leadingZeros_T_189 = _weightQ8_63_5_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_5_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_5_leadingZeros = _weightQ8_63_5_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_5_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_5_expRaw_T_1 = 6'h1f - weightQ8_63_5_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_5_expRaw = weightQ8_63_5_isZero ? 6'h0 : _weightQ8_63_5_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_5_shiftAmt_T_2 = weightQ8_63_5_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_5_shiftAmt = weightQ8_63_5_expRaw > 6'h3 ? _weightQ8_63_5_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_5_mantissaRaw_T = weightQ8_63_5_absClipped >> weightQ8_63_5_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_5_mantissaRaw = _weightQ8_63_5_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_5_mantissa = weightQ8_63_5_expRaw >= 6'h3 ? weightQ8_63_5_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_5_expAdjusted = weightQ8_63_5_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_5_exp_T_4 = weightQ8_63_5_expAdjusted > 7'hf ? 4'hf : weightQ8_63_5_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_5_exp = weightQ8_63_5_isZero ? 4'h0 : _weightQ8_63_5_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_5_fp8 = {weightQ8_63_5_clippedX[31],weightQ8_63_5_exp,weightQ8_63_5_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_6_T = {24'h0,linear_weight_63_6}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_6_sign = _weightQ8_63_6_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_6_absX_T = ~_weightQ8_63_6_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_6_absX_T_2 = _weightQ8_63_6_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_6_absX = weightQ8_63_6_sign ? _weightQ8_63_6_absX_T_2 : _weightQ8_63_6_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_6_shiftedX_T_1 = _GEN_14432 - weightQ8_63_6_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_6_shiftedX_T_3 = weightQ8_63_6_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_6_shiftedX = weightQ8_63_6_sign ? _weightQ8_63_6_shiftedX_T_1 : _weightQ8_63_6_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_6_scaledX_T_1 = weightQ8_63_6_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_6_scaledX = _weightQ8_63_6_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_6_clippedX_T_2 = weightQ8_63_6_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_6_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_6_clippedX = weightQ8_63_6_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_6_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_6_absClipped_T_1 = ~weightQ8_63_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_6_absClipped_T_3 = _weightQ8_63_6_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_6_absClipped = weightQ8_63_6_clippedX[31] ? _weightQ8_63_6_absClipped_T_3 :
    weightQ8_63_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_6_isZero = weightQ8_63_6_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37380 = {{16'd0}, weightQ8_63_6_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_4 = _GEN_37380 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_6 = {weightQ8_63_6_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_8 = _weightQ8_63_6_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_9 = _weightQ8_63_6_leadingZeros_T_4 | _weightQ8_63_6_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37381 = {{8'd0}, _weightQ8_63_6_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_14 = _GEN_37381 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_16 = {_weightQ8_63_6_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_18 = _weightQ8_63_6_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_19 = _weightQ8_63_6_leadingZeros_T_14 | _weightQ8_63_6_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37382 = {{4'd0}, _weightQ8_63_6_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_24 = _GEN_37382 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_26 = {_weightQ8_63_6_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_28 = _weightQ8_63_6_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_29 = _weightQ8_63_6_leadingZeros_T_24 | _weightQ8_63_6_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37383 = {{2'd0}, _weightQ8_63_6_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_34 = _GEN_37383 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_36 = {_weightQ8_63_6_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_38 = _weightQ8_63_6_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_39 = _weightQ8_63_6_leadingZeros_T_34 | _weightQ8_63_6_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37384 = {{1'd0}, _weightQ8_63_6_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_44 = _GEN_37384 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_46 = {_weightQ8_63_6_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_48 = _weightQ8_63_6_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_6_leadingZeros_T_49 = _weightQ8_63_6_leadingZeros_T_44 | _weightQ8_63_6_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37385 = {{8'd0}, weightQ8_63_6_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_55 = _GEN_37385 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_57 = {weightQ8_63_6_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_59 = _weightQ8_63_6_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_60 = _weightQ8_63_6_leadingZeros_T_55 | _weightQ8_63_6_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37386 = {{4'd0}, _weightQ8_63_6_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_65 = _GEN_37386 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_67 = {_weightQ8_63_6_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_69 = _weightQ8_63_6_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_70 = _weightQ8_63_6_leadingZeros_T_65 | _weightQ8_63_6_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37387 = {{2'd0}, _weightQ8_63_6_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_75 = _GEN_37387 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_77 = {_weightQ8_63_6_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_79 = _weightQ8_63_6_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_80 = _weightQ8_63_6_leadingZeros_T_75 | _weightQ8_63_6_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37388 = {{1'd0}, _weightQ8_63_6_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_85 = _GEN_37388 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_87 = {_weightQ8_63_6_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_89 = _weightQ8_63_6_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_6_leadingZeros_T_90 = _weightQ8_63_6_leadingZeros_T_85 | _weightQ8_63_6_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_6_leadingZeros_T_93 = {_weightQ8_63_6_leadingZeros_T_49,_weightQ8_63_6_leadingZeros_T_90,
    weightQ8_63_6_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_143 = _weightQ8_63_6_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_144 = _weightQ8_63_6_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_6_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_145 = _weightQ8_63_6_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_6_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_146 = _weightQ8_63_6_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_6_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_147 = _weightQ8_63_6_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_6_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_148 = _weightQ8_63_6_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_6_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_149 = _weightQ8_63_6_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_6_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_150 = _weightQ8_63_6_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_6_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_151 = _weightQ8_63_6_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_6_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_152 = _weightQ8_63_6_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_6_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_153 = _weightQ8_63_6_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_6_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_154 = _weightQ8_63_6_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_6_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_155 = _weightQ8_63_6_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_6_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_156 = _weightQ8_63_6_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_6_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_157 = _weightQ8_63_6_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_6_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_158 = _weightQ8_63_6_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_6_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_159 = _weightQ8_63_6_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_6_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_160 = _weightQ8_63_6_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_6_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_161 = _weightQ8_63_6_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_6_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_162 = _weightQ8_63_6_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_6_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_163 = _weightQ8_63_6_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_6_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_164 = _weightQ8_63_6_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_6_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_165 = _weightQ8_63_6_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_6_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_166 = _weightQ8_63_6_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_6_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_167 = _weightQ8_63_6_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_6_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_168 = _weightQ8_63_6_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_6_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_169 = _weightQ8_63_6_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_6_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_170 = _weightQ8_63_6_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_6_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_171 = _weightQ8_63_6_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_6_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_172 = _weightQ8_63_6_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_6_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_173 = _weightQ8_63_6_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_6_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_174 = _weightQ8_63_6_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_6_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_175 = _weightQ8_63_6_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_6_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_176 = _weightQ8_63_6_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_6_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_177 = _weightQ8_63_6_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_6_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_178 = _weightQ8_63_6_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_6_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_179 = _weightQ8_63_6_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_6_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_180 = _weightQ8_63_6_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_6_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_181 = _weightQ8_63_6_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_6_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_182 = _weightQ8_63_6_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_6_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_183 = _weightQ8_63_6_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_6_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_184 = _weightQ8_63_6_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_6_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_185 = _weightQ8_63_6_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_6_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_186 = _weightQ8_63_6_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_6_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_187 = _weightQ8_63_6_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_6_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_188 = _weightQ8_63_6_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_6_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_leadingZeros_T_189 = _weightQ8_63_6_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_6_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_6_leadingZeros = _weightQ8_63_6_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_6_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_6_expRaw_T_1 = 6'h1f - weightQ8_63_6_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_6_expRaw = weightQ8_63_6_isZero ? 6'h0 : _weightQ8_63_6_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_6_shiftAmt_T_2 = weightQ8_63_6_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_6_shiftAmt = weightQ8_63_6_expRaw > 6'h3 ? _weightQ8_63_6_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_6_mantissaRaw_T = weightQ8_63_6_absClipped >> weightQ8_63_6_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_6_mantissaRaw = _weightQ8_63_6_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_6_mantissa = weightQ8_63_6_expRaw >= 6'h3 ? weightQ8_63_6_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_6_expAdjusted = weightQ8_63_6_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_6_exp_T_4 = weightQ8_63_6_expAdjusted > 7'hf ? 4'hf : weightQ8_63_6_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_6_exp = weightQ8_63_6_isZero ? 4'h0 : _weightQ8_63_6_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_6_fp8 = {weightQ8_63_6_clippedX[31],weightQ8_63_6_exp,weightQ8_63_6_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_7_T = {24'h0,linear_weight_63_7}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_7_sign = _weightQ8_63_7_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_7_absX_T = ~_weightQ8_63_7_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_7_absX_T_2 = _weightQ8_63_7_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_7_absX = weightQ8_63_7_sign ? _weightQ8_63_7_absX_T_2 : _weightQ8_63_7_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_7_shiftedX_T_1 = _GEN_14432 - weightQ8_63_7_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_7_shiftedX_T_3 = weightQ8_63_7_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_7_shiftedX = weightQ8_63_7_sign ? _weightQ8_63_7_shiftedX_T_1 : _weightQ8_63_7_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_7_scaledX_T_1 = weightQ8_63_7_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_7_scaledX = _weightQ8_63_7_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_7_clippedX_T_2 = weightQ8_63_7_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_7_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_7_clippedX = weightQ8_63_7_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_7_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_7_absClipped_T_1 = ~weightQ8_63_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_7_absClipped_T_3 = _weightQ8_63_7_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_7_absClipped = weightQ8_63_7_clippedX[31] ? _weightQ8_63_7_absClipped_T_3 :
    weightQ8_63_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_7_isZero = weightQ8_63_7_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37391 = {{16'd0}, weightQ8_63_7_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_4 = _GEN_37391 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_6 = {weightQ8_63_7_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_8 = _weightQ8_63_7_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_9 = _weightQ8_63_7_leadingZeros_T_4 | _weightQ8_63_7_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37392 = {{8'd0}, _weightQ8_63_7_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_14 = _GEN_37392 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_16 = {_weightQ8_63_7_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_18 = _weightQ8_63_7_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_19 = _weightQ8_63_7_leadingZeros_T_14 | _weightQ8_63_7_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37393 = {{4'd0}, _weightQ8_63_7_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_24 = _GEN_37393 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_26 = {_weightQ8_63_7_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_28 = _weightQ8_63_7_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_29 = _weightQ8_63_7_leadingZeros_T_24 | _weightQ8_63_7_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37394 = {{2'd0}, _weightQ8_63_7_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_34 = _GEN_37394 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_36 = {_weightQ8_63_7_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_38 = _weightQ8_63_7_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_39 = _weightQ8_63_7_leadingZeros_T_34 | _weightQ8_63_7_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37395 = {{1'd0}, _weightQ8_63_7_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_44 = _GEN_37395 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_46 = {_weightQ8_63_7_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_48 = _weightQ8_63_7_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_7_leadingZeros_T_49 = _weightQ8_63_7_leadingZeros_T_44 | _weightQ8_63_7_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37396 = {{8'd0}, weightQ8_63_7_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_55 = _GEN_37396 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_57 = {weightQ8_63_7_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_59 = _weightQ8_63_7_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_60 = _weightQ8_63_7_leadingZeros_T_55 | _weightQ8_63_7_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37397 = {{4'd0}, _weightQ8_63_7_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_65 = _GEN_37397 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_67 = {_weightQ8_63_7_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_69 = _weightQ8_63_7_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_70 = _weightQ8_63_7_leadingZeros_T_65 | _weightQ8_63_7_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37398 = {{2'd0}, _weightQ8_63_7_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_75 = _GEN_37398 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_77 = {_weightQ8_63_7_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_79 = _weightQ8_63_7_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_80 = _weightQ8_63_7_leadingZeros_T_75 | _weightQ8_63_7_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37399 = {{1'd0}, _weightQ8_63_7_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_85 = _GEN_37399 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_87 = {_weightQ8_63_7_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_89 = _weightQ8_63_7_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_7_leadingZeros_T_90 = _weightQ8_63_7_leadingZeros_T_85 | _weightQ8_63_7_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_7_leadingZeros_T_93 = {_weightQ8_63_7_leadingZeros_T_49,_weightQ8_63_7_leadingZeros_T_90,
    weightQ8_63_7_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_143 = _weightQ8_63_7_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_144 = _weightQ8_63_7_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_7_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_145 = _weightQ8_63_7_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_7_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_146 = _weightQ8_63_7_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_7_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_147 = _weightQ8_63_7_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_7_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_148 = _weightQ8_63_7_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_7_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_149 = _weightQ8_63_7_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_7_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_150 = _weightQ8_63_7_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_7_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_151 = _weightQ8_63_7_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_7_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_152 = _weightQ8_63_7_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_7_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_153 = _weightQ8_63_7_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_7_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_154 = _weightQ8_63_7_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_7_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_155 = _weightQ8_63_7_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_7_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_156 = _weightQ8_63_7_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_7_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_157 = _weightQ8_63_7_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_7_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_158 = _weightQ8_63_7_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_7_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_159 = _weightQ8_63_7_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_7_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_160 = _weightQ8_63_7_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_7_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_161 = _weightQ8_63_7_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_7_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_162 = _weightQ8_63_7_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_7_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_163 = _weightQ8_63_7_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_7_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_164 = _weightQ8_63_7_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_7_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_165 = _weightQ8_63_7_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_7_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_166 = _weightQ8_63_7_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_7_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_167 = _weightQ8_63_7_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_7_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_168 = _weightQ8_63_7_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_7_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_169 = _weightQ8_63_7_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_7_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_170 = _weightQ8_63_7_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_7_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_171 = _weightQ8_63_7_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_7_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_172 = _weightQ8_63_7_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_7_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_173 = _weightQ8_63_7_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_7_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_174 = _weightQ8_63_7_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_7_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_175 = _weightQ8_63_7_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_7_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_176 = _weightQ8_63_7_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_7_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_177 = _weightQ8_63_7_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_7_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_178 = _weightQ8_63_7_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_7_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_179 = _weightQ8_63_7_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_7_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_180 = _weightQ8_63_7_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_7_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_181 = _weightQ8_63_7_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_7_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_182 = _weightQ8_63_7_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_7_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_183 = _weightQ8_63_7_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_7_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_184 = _weightQ8_63_7_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_7_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_185 = _weightQ8_63_7_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_7_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_186 = _weightQ8_63_7_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_7_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_187 = _weightQ8_63_7_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_7_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_188 = _weightQ8_63_7_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_7_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_leadingZeros_T_189 = _weightQ8_63_7_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_7_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_7_leadingZeros = _weightQ8_63_7_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_7_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_7_expRaw_T_1 = 6'h1f - weightQ8_63_7_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_7_expRaw = weightQ8_63_7_isZero ? 6'h0 : _weightQ8_63_7_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_7_shiftAmt_T_2 = weightQ8_63_7_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_7_shiftAmt = weightQ8_63_7_expRaw > 6'h3 ? _weightQ8_63_7_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_7_mantissaRaw_T = weightQ8_63_7_absClipped >> weightQ8_63_7_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_7_mantissaRaw = _weightQ8_63_7_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_7_mantissa = weightQ8_63_7_expRaw >= 6'h3 ? weightQ8_63_7_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_7_expAdjusted = weightQ8_63_7_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_7_exp_T_4 = weightQ8_63_7_expAdjusted > 7'hf ? 4'hf : weightQ8_63_7_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_7_exp = weightQ8_63_7_isZero ? 4'h0 : _weightQ8_63_7_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_7_fp8 = {weightQ8_63_7_clippedX[31],weightQ8_63_7_exp,weightQ8_63_7_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_8_T = {24'h0,linear_weight_63_8}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_8_sign = _weightQ8_63_8_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_8_absX_T = ~_weightQ8_63_8_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_8_absX_T_2 = _weightQ8_63_8_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_8_absX = weightQ8_63_8_sign ? _weightQ8_63_8_absX_T_2 : _weightQ8_63_8_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_8_shiftedX_T_1 = _GEN_14432 - weightQ8_63_8_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_8_shiftedX_T_3 = weightQ8_63_8_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_8_shiftedX = weightQ8_63_8_sign ? _weightQ8_63_8_shiftedX_T_1 : _weightQ8_63_8_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_8_scaledX_T_1 = weightQ8_63_8_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_8_scaledX = _weightQ8_63_8_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_8_clippedX_T_2 = weightQ8_63_8_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_8_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_8_clippedX = weightQ8_63_8_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_8_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_8_absClipped_T_1 = ~weightQ8_63_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_8_absClipped_T_3 = _weightQ8_63_8_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_8_absClipped = weightQ8_63_8_clippedX[31] ? _weightQ8_63_8_absClipped_T_3 :
    weightQ8_63_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_8_isZero = weightQ8_63_8_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37402 = {{16'd0}, weightQ8_63_8_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_4 = _GEN_37402 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_6 = {weightQ8_63_8_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_8 = _weightQ8_63_8_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_9 = _weightQ8_63_8_leadingZeros_T_4 | _weightQ8_63_8_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37403 = {{8'd0}, _weightQ8_63_8_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_14 = _GEN_37403 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_16 = {_weightQ8_63_8_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_18 = _weightQ8_63_8_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_19 = _weightQ8_63_8_leadingZeros_T_14 | _weightQ8_63_8_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37404 = {{4'd0}, _weightQ8_63_8_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_24 = _GEN_37404 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_26 = {_weightQ8_63_8_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_28 = _weightQ8_63_8_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_29 = _weightQ8_63_8_leadingZeros_T_24 | _weightQ8_63_8_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37405 = {{2'd0}, _weightQ8_63_8_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_34 = _GEN_37405 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_36 = {_weightQ8_63_8_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_38 = _weightQ8_63_8_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_39 = _weightQ8_63_8_leadingZeros_T_34 | _weightQ8_63_8_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37406 = {{1'd0}, _weightQ8_63_8_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_44 = _GEN_37406 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_46 = {_weightQ8_63_8_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_48 = _weightQ8_63_8_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_8_leadingZeros_T_49 = _weightQ8_63_8_leadingZeros_T_44 | _weightQ8_63_8_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37407 = {{8'd0}, weightQ8_63_8_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_55 = _GEN_37407 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_57 = {weightQ8_63_8_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_59 = _weightQ8_63_8_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_60 = _weightQ8_63_8_leadingZeros_T_55 | _weightQ8_63_8_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37408 = {{4'd0}, _weightQ8_63_8_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_65 = _GEN_37408 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_67 = {_weightQ8_63_8_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_69 = _weightQ8_63_8_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_70 = _weightQ8_63_8_leadingZeros_T_65 | _weightQ8_63_8_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37409 = {{2'd0}, _weightQ8_63_8_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_75 = _GEN_37409 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_77 = {_weightQ8_63_8_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_79 = _weightQ8_63_8_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_80 = _weightQ8_63_8_leadingZeros_T_75 | _weightQ8_63_8_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37410 = {{1'd0}, _weightQ8_63_8_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_85 = _GEN_37410 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_87 = {_weightQ8_63_8_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_89 = _weightQ8_63_8_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_8_leadingZeros_T_90 = _weightQ8_63_8_leadingZeros_T_85 | _weightQ8_63_8_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_8_leadingZeros_T_93 = {_weightQ8_63_8_leadingZeros_T_49,_weightQ8_63_8_leadingZeros_T_90,
    weightQ8_63_8_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_143 = _weightQ8_63_8_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_144 = _weightQ8_63_8_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_8_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_145 = _weightQ8_63_8_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_8_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_146 = _weightQ8_63_8_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_8_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_147 = _weightQ8_63_8_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_8_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_148 = _weightQ8_63_8_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_8_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_149 = _weightQ8_63_8_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_8_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_150 = _weightQ8_63_8_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_8_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_151 = _weightQ8_63_8_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_8_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_152 = _weightQ8_63_8_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_8_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_153 = _weightQ8_63_8_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_8_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_154 = _weightQ8_63_8_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_8_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_155 = _weightQ8_63_8_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_8_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_156 = _weightQ8_63_8_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_8_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_157 = _weightQ8_63_8_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_8_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_158 = _weightQ8_63_8_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_8_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_159 = _weightQ8_63_8_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_8_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_160 = _weightQ8_63_8_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_8_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_161 = _weightQ8_63_8_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_8_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_162 = _weightQ8_63_8_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_8_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_163 = _weightQ8_63_8_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_8_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_164 = _weightQ8_63_8_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_8_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_165 = _weightQ8_63_8_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_8_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_166 = _weightQ8_63_8_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_8_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_167 = _weightQ8_63_8_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_8_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_168 = _weightQ8_63_8_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_8_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_169 = _weightQ8_63_8_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_8_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_170 = _weightQ8_63_8_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_8_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_171 = _weightQ8_63_8_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_8_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_172 = _weightQ8_63_8_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_8_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_173 = _weightQ8_63_8_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_8_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_174 = _weightQ8_63_8_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_8_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_175 = _weightQ8_63_8_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_8_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_176 = _weightQ8_63_8_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_8_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_177 = _weightQ8_63_8_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_8_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_178 = _weightQ8_63_8_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_8_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_179 = _weightQ8_63_8_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_8_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_180 = _weightQ8_63_8_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_8_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_181 = _weightQ8_63_8_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_8_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_182 = _weightQ8_63_8_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_8_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_183 = _weightQ8_63_8_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_8_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_184 = _weightQ8_63_8_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_8_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_185 = _weightQ8_63_8_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_8_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_186 = _weightQ8_63_8_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_8_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_187 = _weightQ8_63_8_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_8_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_188 = _weightQ8_63_8_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_8_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_leadingZeros_T_189 = _weightQ8_63_8_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_8_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_8_leadingZeros = _weightQ8_63_8_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_8_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_8_expRaw_T_1 = 6'h1f - weightQ8_63_8_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_8_expRaw = weightQ8_63_8_isZero ? 6'h0 : _weightQ8_63_8_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_8_shiftAmt_T_2 = weightQ8_63_8_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_8_shiftAmt = weightQ8_63_8_expRaw > 6'h3 ? _weightQ8_63_8_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_8_mantissaRaw_T = weightQ8_63_8_absClipped >> weightQ8_63_8_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_8_mantissaRaw = _weightQ8_63_8_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_8_mantissa = weightQ8_63_8_expRaw >= 6'h3 ? weightQ8_63_8_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_8_expAdjusted = weightQ8_63_8_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_8_exp_T_4 = weightQ8_63_8_expAdjusted > 7'hf ? 4'hf : weightQ8_63_8_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_8_exp = weightQ8_63_8_isZero ? 4'h0 : _weightQ8_63_8_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_8_fp8 = {weightQ8_63_8_clippedX[31],weightQ8_63_8_exp,weightQ8_63_8_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_9_T = {24'h0,linear_weight_63_9}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_9_sign = _weightQ8_63_9_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_9_absX_T = ~_weightQ8_63_9_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_9_absX_T_2 = _weightQ8_63_9_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_9_absX = weightQ8_63_9_sign ? _weightQ8_63_9_absX_T_2 : _weightQ8_63_9_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_9_shiftedX_T_1 = _GEN_14432 - weightQ8_63_9_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_9_shiftedX_T_3 = weightQ8_63_9_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_9_shiftedX = weightQ8_63_9_sign ? _weightQ8_63_9_shiftedX_T_1 : _weightQ8_63_9_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_9_scaledX_T_1 = weightQ8_63_9_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_9_scaledX = _weightQ8_63_9_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_9_clippedX_T_2 = weightQ8_63_9_scaledX < 49'hfffffe40 ? 49'hfffffe40 : weightQ8_63_9_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_9_clippedX = weightQ8_63_9_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_9_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_9_absClipped_T_1 = ~weightQ8_63_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_9_absClipped_T_3 = _weightQ8_63_9_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_9_absClipped = weightQ8_63_9_clippedX[31] ? _weightQ8_63_9_absClipped_T_3 :
    weightQ8_63_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_9_isZero = weightQ8_63_9_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37413 = {{16'd0}, weightQ8_63_9_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_4 = _GEN_37413 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_6 = {weightQ8_63_9_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_8 = _weightQ8_63_9_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_9 = _weightQ8_63_9_leadingZeros_T_4 | _weightQ8_63_9_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37414 = {{8'd0}, _weightQ8_63_9_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_14 = _GEN_37414 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_16 = {_weightQ8_63_9_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_18 = _weightQ8_63_9_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_19 = _weightQ8_63_9_leadingZeros_T_14 | _weightQ8_63_9_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37415 = {{4'd0}, _weightQ8_63_9_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_24 = _GEN_37415 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_26 = {_weightQ8_63_9_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_28 = _weightQ8_63_9_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_29 = _weightQ8_63_9_leadingZeros_T_24 | _weightQ8_63_9_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37416 = {{2'd0}, _weightQ8_63_9_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_34 = _GEN_37416 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_36 = {_weightQ8_63_9_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_38 = _weightQ8_63_9_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_39 = _weightQ8_63_9_leadingZeros_T_34 | _weightQ8_63_9_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37417 = {{1'd0}, _weightQ8_63_9_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_44 = _GEN_37417 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_46 = {_weightQ8_63_9_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_48 = _weightQ8_63_9_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_9_leadingZeros_T_49 = _weightQ8_63_9_leadingZeros_T_44 | _weightQ8_63_9_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37418 = {{8'd0}, weightQ8_63_9_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_55 = _GEN_37418 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_57 = {weightQ8_63_9_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_59 = _weightQ8_63_9_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_60 = _weightQ8_63_9_leadingZeros_T_55 | _weightQ8_63_9_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37419 = {{4'd0}, _weightQ8_63_9_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_65 = _GEN_37419 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_67 = {_weightQ8_63_9_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_69 = _weightQ8_63_9_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_70 = _weightQ8_63_9_leadingZeros_T_65 | _weightQ8_63_9_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37420 = {{2'd0}, _weightQ8_63_9_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_75 = _GEN_37420 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_77 = {_weightQ8_63_9_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_79 = _weightQ8_63_9_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_80 = _weightQ8_63_9_leadingZeros_T_75 | _weightQ8_63_9_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37421 = {{1'd0}, _weightQ8_63_9_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_85 = _GEN_37421 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_87 = {_weightQ8_63_9_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_89 = _weightQ8_63_9_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_9_leadingZeros_T_90 = _weightQ8_63_9_leadingZeros_T_85 | _weightQ8_63_9_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_9_leadingZeros_T_93 = {_weightQ8_63_9_leadingZeros_T_49,_weightQ8_63_9_leadingZeros_T_90,
    weightQ8_63_9_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_143 = _weightQ8_63_9_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_144 = _weightQ8_63_9_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_9_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_145 = _weightQ8_63_9_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_9_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_146 = _weightQ8_63_9_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_9_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_147 = _weightQ8_63_9_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_9_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_148 = _weightQ8_63_9_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_9_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_149 = _weightQ8_63_9_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_9_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_150 = _weightQ8_63_9_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_9_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_151 = _weightQ8_63_9_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_9_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_152 = _weightQ8_63_9_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_9_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_153 = _weightQ8_63_9_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_9_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_154 = _weightQ8_63_9_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_9_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_155 = _weightQ8_63_9_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_9_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_156 = _weightQ8_63_9_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_9_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_157 = _weightQ8_63_9_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_9_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_158 = _weightQ8_63_9_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_9_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_159 = _weightQ8_63_9_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_9_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_160 = _weightQ8_63_9_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_9_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_161 = _weightQ8_63_9_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_9_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_162 = _weightQ8_63_9_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_9_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_163 = _weightQ8_63_9_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_9_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_164 = _weightQ8_63_9_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_9_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_165 = _weightQ8_63_9_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_9_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_166 = _weightQ8_63_9_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_9_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_167 = _weightQ8_63_9_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_9_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_168 = _weightQ8_63_9_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_9_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_169 = _weightQ8_63_9_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_9_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_170 = _weightQ8_63_9_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_9_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_171 = _weightQ8_63_9_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_9_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_172 = _weightQ8_63_9_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_9_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_173 = _weightQ8_63_9_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_9_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_174 = _weightQ8_63_9_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_9_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_175 = _weightQ8_63_9_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_9_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_176 = _weightQ8_63_9_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_9_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_177 = _weightQ8_63_9_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_9_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_178 = _weightQ8_63_9_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_9_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_179 = _weightQ8_63_9_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_9_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_180 = _weightQ8_63_9_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_9_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_181 = _weightQ8_63_9_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_9_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_182 = _weightQ8_63_9_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_9_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_183 = _weightQ8_63_9_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_9_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_184 = _weightQ8_63_9_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_9_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_185 = _weightQ8_63_9_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_9_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_186 = _weightQ8_63_9_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_9_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_187 = _weightQ8_63_9_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_9_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_188 = _weightQ8_63_9_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_9_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_leadingZeros_T_189 = _weightQ8_63_9_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_9_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_9_leadingZeros = _weightQ8_63_9_leadingZeros_T_93[0] ? 6'h0 : _weightQ8_63_9_leadingZeros_T_189
    ; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_9_expRaw_T_1 = 6'h1f - weightQ8_63_9_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_9_expRaw = weightQ8_63_9_isZero ? 6'h0 : _weightQ8_63_9_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_9_shiftAmt_T_2 = weightQ8_63_9_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_9_shiftAmt = weightQ8_63_9_expRaw > 6'h3 ? _weightQ8_63_9_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_9_mantissaRaw_T = weightQ8_63_9_absClipped >> weightQ8_63_9_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_9_mantissaRaw = _weightQ8_63_9_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_9_mantissa = weightQ8_63_9_expRaw >= 6'h3 ? weightQ8_63_9_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_9_expAdjusted = weightQ8_63_9_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_9_exp_T_4 = weightQ8_63_9_expAdjusted > 7'hf ? 4'hf : weightQ8_63_9_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_9_exp = weightQ8_63_9_isZero ? 4'h0 : _weightQ8_63_9_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_9_fp8 = {weightQ8_63_9_clippedX[31],weightQ8_63_9_exp,weightQ8_63_9_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_10_T = {24'h0,linear_weight_63_10}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_10_sign = _weightQ8_63_10_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_10_absX_T = ~_weightQ8_63_10_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_10_absX_T_2 = _weightQ8_63_10_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_10_absX = weightQ8_63_10_sign ? _weightQ8_63_10_absX_T_2 : _weightQ8_63_10_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_10_shiftedX_T_1 = _GEN_14432 - weightQ8_63_10_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_10_shiftedX_T_3 = weightQ8_63_10_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_10_shiftedX = weightQ8_63_10_sign ? _weightQ8_63_10_shiftedX_T_1 :
    _weightQ8_63_10_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_10_scaledX_T_1 = weightQ8_63_10_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_10_scaledX = _weightQ8_63_10_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_10_clippedX_T_2 = weightQ8_63_10_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_10_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_10_clippedX = weightQ8_63_10_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_10_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_10_absClipped_T_1 = ~weightQ8_63_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_10_absClipped_T_3 = _weightQ8_63_10_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_10_absClipped = weightQ8_63_10_clippedX[31] ? _weightQ8_63_10_absClipped_T_3 :
    weightQ8_63_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_10_isZero = weightQ8_63_10_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37424 = {{16'd0}, weightQ8_63_10_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_4 = _GEN_37424 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_6 = {weightQ8_63_10_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_8 = _weightQ8_63_10_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_9 = _weightQ8_63_10_leadingZeros_T_4 | _weightQ8_63_10_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37425 = {{8'd0}, _weightQ8_63_10_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_14 = _GEN_37425 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_16 = {_weightQ8_63_10_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_18 = _weightQ8_63_10_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_19 = _weightQ8_63_10_leadingZeros_T_14 | _weightQ8_63_10_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37426 = {{4'd0}, _weightQ8_63_10_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_24 = _GEN_37426 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_26 = {_weightQ8_63_10_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_28 = _weightQ8_63_10_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_29 = _weightQ8_63_10_leadingZeros_T_24 | _weightQ8_63_10_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37427 = {{2'd0}, _weightQ8_63_10_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_34 = _GEN_37427 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_36 = {_weightQ8_63_10_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_38 = _weightQ8_63_10_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_39 = _weightQ8_63_10_leadingZeros_T_34 | _weightQ8_63_10_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37428 = {{1'd0}, _weightQ8_63_10_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_44 = _GEN_37428 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_46 = {_weightQ8_63_10_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_48 = _weightQ8_63_10_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_10_leadingZeros_T_49 = _weightQ8_63_10_leadingZeros_T_44 | _weightQ8_63_10_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37429 = {{8'd0}, weightQ8_63_10_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_55 = _GEN_37429 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_57 = {weightQ8_63_10_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_59 = _weightQ8_63_10_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_60 = _weightQ8_63_10_leadingZeros_T_55 | _weightQ8_63_10_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37430 = {{4'd0}, _weightQ8_63_10_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_65 = _GEN_37430 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_67 = {_weightQ8_63_10_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_69 = _weightQ8_63_10_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_70 = _weightQ8_63_10_leadingZeros_T_65 | _weightQ8_63_10_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37431 = {{2'd0}, _weightQ8_63_10_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_75 = _GEN_37431 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_77 = {_weightQ8_63_10_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_79 = _weightQ8_63_10_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_80 = _weightQ8_63_10_leadingZeros_T_75 | _weightQ8_63_10_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37432 = {{1'd0}, _weightQ8_63_10_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_85 = _GEN_37432 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_87 = {_weightQ8_63_10_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_89 = _weightQ8_63_10_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_10_leadingZeros_T_90 = _weightQ8_63_10_leadingZeros_T_85 | _weightQ8_63_10_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_10_leadingZeros_T_93 = {_weightQ8_63_10_leadingZeros_T_49,_weightQ8_63_10_leadingZeros_T_90,
    weightQ8_63_10_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_143 = _weightQ8_63_10_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_144 = _weightQ8_63_10_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_10_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_145 = _weightQ8_63_10_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_10_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_146 = _weightQ8_63_10_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_10_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_147 = _weightQ8_63_10_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_10_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_148 = _weightQ8_63_10_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_10_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_149 = _weightQ8_63_10_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_10_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_150 = _weightQ8_63_10_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_10_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_151 = _weightQ8_63_10_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_10_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_152 = _weightQ8_63_10_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_10_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_153 = _weightQ8_63_10_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_10_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_154 = _weightQ8_63_10_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_10_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_155 = _weightQ8_63_10_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_10_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_156 = _weightQ8_63_10_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_10_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_157 = _weightQ8_63_10_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_10_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_158 = _weightQ8_63_10_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_10_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_159 = _weightQ8_63_10_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_10_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_160 = _weightQ8_63_10_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_10_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_161 = _weightQ8_63_10_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_10_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_162 = _weightQ8_63_10_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_10_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_163 = _weightQ8_63_10_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_10_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_164 = _weightQ8_63_10_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_10_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_165 = _weightQ8_63_10_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_10_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_166 = _weightQ8_63_10_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_10_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_167 = _weightQ8_63_10_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_10_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_168 = _weightQ8_63_10_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_10_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_169 = _weightQ8_63_10_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_10_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_170 = _weightQ8_63_10_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_10_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_171 = _weightQ8_63_10_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_10_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_172 = _weightQ8_63_10_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_10_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_173 = _weightQ8_63_10_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_10_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_174 = _weightQ8_63_10_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_10_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_175 = _weightQ8_63_10_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_10_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_176 = _weightQ8_63_10_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_10_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_177 = _weightQ8_63_10_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_10_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_178 = _weightQ8_63_10_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_10_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_179 = _weightQ8_63_10_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_10_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_180 = _weightQ8_63_10_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_10_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_181 = _weightQ8_63_10_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_10_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_182 = _weightQ8_63_10_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_10_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_183 = _weightQ8_63_10_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_10_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_184 = _weightQ8_63_10_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_10_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_185 = _weightQ8_63_10_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_10_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_186 = _weightQ8_63_10_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_10_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_187 = _weightQ8_63_10_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_10_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_188 = _weightQ8_63_10_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_10_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_leadingZeros_T_189 = _weightQ8_63_10_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_10_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_10_leadingZeros = _weightQ8_63_10_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_10_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_10_expRaw_T_1 = 6'h1f - weightQ8_63_10_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_10_expRaw = weightQ8_63_10_isZero ? 6'h0 : _weightQ8_63_10_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_10_shiftAmt_T_2 = weightQ8_63_10_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_10_shiftAmt = weightQ8_63_10_expRaw > 6'h3 ? _weightQ8_63_10_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_10_mantissaRaw_T = weightQ8_63_10_absClipped >> weightQ8_63_10_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_10_mantissaRaw = _weightQ8_63_10_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_10_mantissa = weightQ8_63_10_expRaw >= 6'h3 ? weightQ8_63_10_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_10_expAdjusted = weightQ8_63_10_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_10_exp_T_4 = weightQ8_63_10_expAdjusted > 7'hf ? 4'hf : weightQ8_63_10_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_10_exp = weightQ8_63_10_isZero ? 4'h0 : _weightQ8_63_10_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_10_fp8 = {weightQ8_63_10_clippedX[31],weightQ8_63_10_exp,weightQ8_63_10_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_11_T = {24'h0,linear_weight_63_11}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_11_sign = _weightQ8_63_11_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_11_absX_T = ~_weightQ8_63_11_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_11_absX_T_2 = _weightQ8_63_11_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_11_absX = weightQ8_63_11_sign ? _weightQ8_63_11_absX_T_2 : _weightQ8_63_11_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_11_shiftedX_T_1 = _GEN_14432 - weightQ8_63_11_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_11_shiftedX_T_3 = weightQ8_63_11_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_11_shiftedX = weightQ8_63_11_sign ? _weightQ8_63_11_shiftedX_T_1 :
    _weightQ8_63_11_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_11_scaledX_T_1 = weightQ8_63_11_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_11_scaledX = _weightQ8_63_11_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_11_clippedX_T_2 = weightQ8_63_11_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_11_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_11_clippedX = weightQ8_63_11_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_11_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_11_absClipped_T_1 = ~weightQ8_63_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_11_absClipped_T_3 = _weightQ8_63_11_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_11_absClipped = weightQ8_63_11_clippedX[31] ? _weightQ8_63_11_absClipped_T_3 :
    weightQ8_63_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_11_isZero = weightQ8_63_11_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37435 = {{16'd0}, weightQ8_63_11_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_4 = _GEN_37435 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_6 = {weightQ8_63_11_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_8 = _weightQ8_63_11_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_9 = _weightQ8_63_11_leadingZeros_T_4 | _weightQ8_63_11_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37436 = {{8'd0}, _weightQ8_63_11_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_14 = _GEN_37436 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_16 = {_weightQ8_63_11_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_18 = _weightQ8_63_11_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_19 = _weightQ8_63_11_leadingZeros_T_14 | _weightQ8_63_11_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37437 = {{4'd0}, _weightQ8_63_11_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_24 = _GEN_37437 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_26 = {_weightQ8_63_11_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_28 = _weightQ8_63_11_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_29 = _weightQ8_63_11_leadingZeros_T_24 | _weightQ8_63_11_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37438 = {{2'd0}, _weightQ8_63_11_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_34 = _GEN_37438 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_36 = {_weightQ8_63_11_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_38 = _weightQ8_63_11_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_39 = _weightQ8_63_11_leadingZeros_T_34 | _weightQ8_63_11_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37439 = {{1'd0}, _weightQ8_63_11_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_44 = _GEN_37439 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_46 = {_weightQ8_63_11_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_48 = _weightQ8_63_11_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_11_leadingZeros_T_49 = _weightQ8_63_11_leadingZeros_T_44 | _weightQ8_63_11_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37440 = {{8'd0}, weightQ8_63_11_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_55 = _GEN_37440 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_57 = {weightQ8_63_11_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_59 = _weightQ8_63_11_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_60 = _weightQ8_63_11_leadingZeros_T_55 | _weightQ8_63_11_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37441 = {{4'd0}, _weightQ8_63_11_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_65 = _GEN_37441 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_67 = {_weightQ8_63_11_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_69 = _weightQ8_63_11_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_70 = _weightQ8_63_11_leadingZeros_T_65 | _weightQ8_63_11_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37442 = {{2'd0}, _weightQ8_63_11_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_75 = _GEN_37442 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_77 = {_weightQ8_63_11_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_79 = _weightQ8_63_11_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_80 = _weightQ8_63_11_leadingZeros_T_75 | _weightQ8_63_11_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37443 = {{1'd0}, _weightQ8_63_11_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_85 = _GEN_37443 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_87 = {_weightQ8_63_11_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_89 = _weightQ8_63_11_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_11_leadingZeros_T_90 = _weightQ8_63_11_leadingZeros_T_85 | _weightQ8_63_11_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_11_leadingZeros_T_93 = {_weightQ8_63_11_leadingZeros_T_49,_weightQ8_63_11_leadingZeros_T_90,
    weightQ8_63_11_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_143 = _weightQ8_63_11_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_144 = _weightQ8_63_11_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_11_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_145 = _weightQ8_63_11_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_11_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_146 = _weightQ8_63_11_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_11_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_147 = _weightQ8_63_11_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_11_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_148 = _weightQ8_63_11_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_11_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_149 = _weightQ8_63_11_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_11_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_150 = _weightQ8_63_11_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_11_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_151 = _weightQ8_63_11_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_11_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_152 = _weightQ8_63_11_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_11_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_153 = _weightQ8_63_11_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_11_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_154 = _weightQ8_63_11_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_11_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_155 = _weightQ8_63_11_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_11_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_156 = _weightQ8_63_11_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_11_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_157 = _weightQ8_63_11_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_11_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_158 = _weightQ8_63_11_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_11_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_159 = _weightQ8_63_11_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_11_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_160 = _weightQ8_63_11_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_11_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_161 = _weightQ8_63_11_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_11_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_162 = _weightQ8_63_11_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_11_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_163 = _weightQ8_63_11_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_11_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_164 = _weightQ8_63_11_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_11_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_165 = _weightQ8_63_11_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_11_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_166 = _weightQ8_63_11_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_11_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_167 = _weightQ8_63_11_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_11_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_168 = _weightQ8_63_11_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_11_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_169 = _weightQ8_63_11_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_11_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_170 = _weightQ8_63_11_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_11_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_171 = _weightQ8_63_11_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_11_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_172 = _weightQ8_63_11_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_11_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_173 = _weightQ8_63_11_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_11_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_174 = _weightQ8_63_11_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_11_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_175 = _weightQ8_63_11_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_11_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_176 = _weightQ8_63_11_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_11_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_177 = _weightQ8_63_11_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_11_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_178 = _weightQ8_63_11_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_11_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_179 = _weightQ8_63_11_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_11_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_180 = _weightQ8_63_11_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_11_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_181 = _weightQ8_63_11_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_11_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_182 = _weightQ8_63_11_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_11_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_183 = _weightQ8_63_11_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_11_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_184 = _weightQ8_63_11_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_11_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_185 = _weightQ8_63_11_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_11_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_186 = _weightQ8_63_11_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_11_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_187 = _weightQ8_63_11_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_11_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_188 = _weightQ8_63_11_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_11_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_leadingZeros_T_189 = _weightQ8_63_11_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_11_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_11_leadingZeros = _weightQ8_63_11_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_11_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_11_expRaw_T_1 = 6'h1f - weightQ8_63_11_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_11_expRaw = weightQ8_63_11_isZero ? 6'h0 : _weightQ8_63_11_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_11_shiftAmt_T_2 = weightQ8_63_11_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_11_shiftAmt = weightQ8_63_11_expRaw > 6'h3 ? _weightQ8_63_11_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_11_mantissaRaw_T = weightQ8_63_11_absClipped >> weightQ8_63_11_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_11_mantissaRaw = _weightQ8_63_11_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_11_mantissa = weightQ8_63_11_expRaw >= 6'h3 ? weightQ8_63_11_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_11_expAdjusted = weightQ8_63_11_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_11_exp_T_4 = weightQ8_63_11_expAdjusted > 7'hf ? 4'hf : weightQ8_63_11_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_11_exp = weightQ8_63_11_isZero ? 4'h0 : _weightQ8_63_11_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_11_fp8 = {weightQ8_63_11_clippedX[31],weightQ8_63_11_exp,weightQ8_63_11_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_12_T = {24'h0,linear_weight_63_12}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_12_sign = _weightQ8_63_12_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_12_absX_T = ~_weightQ8_63_12_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_12_absX_T_2 = _weightQ8_63_12_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_12_absX = weightQ8_63_12_sign ? _weightQ8_63_12_absX_T_2 : _weightQ8_63_12_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_12_shiftedX_T_1 = _GEN_14432 - weightQ8_63_12_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_12_shiftedX_T_3 = weightQ8_63_12_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_12_shiftedX = weightQ8_63_12_sign ? _weightQ8_63_12_shiftedX_T_1 :
    _weightQ8_63_12_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_12_scaledX_T_1 = weightQ8_63_12_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_12_scaledX = _weightQ8_63_12_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_12_clippedX_T_2 = weightQ8_63_12_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_12_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_12_clippedX = weightQ8_63_12_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_12_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_12_absClipped_T_1 = ~weightQ8_63_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_12_absClipped_T_3 = _weightQ8_63_12_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_12_absClipped = weightQ8_63_12_clippedX[31] ? _weightQ8_63_12_absClipped_T_3 :
    weightQ8_63_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_12_isZero = weightQ8_63_12_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37446 = {{16'd0}, weightQ8_63_12_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_4 = _GEN_37446 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_6 = {weightQ8_63_12_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_8 = _weightQ8_63_12_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_9 = _weightQ8_63_12_leadingZeros_T_4 | _weightQ8_63_12_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37447 = {{8'd0}, _weightQ8_63_12_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_14 = _GEN_37447 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_16 = {_weightQ8_63_12_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_18 = _weightQ8_63_12_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_19 = _weightQ8_63_12_leadingZeros_T_14 | _weightQ8_63_12_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37448 = {{4'd0}, _weightQ8_63_12_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_24 = _GEN_37448 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_26 = {_weightQ8_63_12_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_28 = _weightQ8_63_12_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_29 = _weightQ8_63_12_leadingZeros_T_24 | _weightQ8_63_12_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37449 = {{2'd0}, _weightQ8_63_12_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_34 = _GEN_37449 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_36 = {_weightQ8_63_12_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_38 = _weightQ8_63_12_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_39 = _weightQ8_63_12_leadingZeros_T_34 | _weightQ8_63_12_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37450 = {{1'd0}, _weightQ8_63_12_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_44 = _GEN_37450 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_46 = {_weightQ8_63_12_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_48 = _weightQ8_63_12_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_12_leadingZeros_T_49 = _weightQ8_63_12_leadingZeros_T_44 | _weightQ8_63_12_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37451 = {{8'd0}, weightQ8_63_12_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_55 = _GEN_37451 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_57 = {weightQ8_63_12_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_59 = _weightQ8_63_12_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_60 = _weightQ8_63_12_leadingZeros_T_55 | _weightQ8_63_12_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37452 = {{4'd0}, _weightQ8_63_12_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_65 = _GEN_37452 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_67 = {_weightQ8_63_12_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_69 = _weightQ8_63_12_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_70 = _weightQ8_63_12_leadingZeros_T_65 | _weightQ8_63_12_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37453 = {{2'd0}, _weightQ8_63_12_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_75 = _GEN_37453 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_77 = {_weightQ8_63_12_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_79 = _weightQ8_63_12_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_80 = _weightQ8_63_12_leadingZeros_T_75 | _weightQ8_63_12_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37454 = {{1'd0}, _weightQ8_63_12_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_85 = _GEN_37454 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_87 = {_weightQ8_63_12_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_89 = _weightQ8_63_12_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_12_leadingZeros_T_90 = _weightQ8_63_12_leadingZeros_T_85 | _weightQ8_63_12_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_12_leadingZeros_T_93 = {_weightQ8_63_12_leadingZeros_T_49,_weightQ8_63_12_leadingZeros_T_90,
    weightQ8_63_12_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_143 = _weightQ8_63_12_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_144 = _weightQ8_63_12_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_12_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_145 = _weightQ8_63_12_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_12_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_146 = _weightQ8_63_12_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_12_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_147 = _weightQ8_63_12_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_12_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_148 = _weightQ8_63_12_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_12_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_149 = _weightQ8_63_12_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_12_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_150 = _weightQ8_63_12_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_12_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_151 = _weightQ8_63_12_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_12_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_152 = _weightQ8_63_12_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_12_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_153 = _weightQ8_63_12_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_12_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_154 = _weightQ8_63_12_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_12_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_155 = _weightQ8_63_12_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_12_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_156 = _weightQ8_63_12_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_12_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_157 = _weightQ8_63_12_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_12_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_158 = _weightQ8_63_12_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_12_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_159 = _weightQ8_63_12_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_12_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_160 = _weightQ8_63_12_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_12_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_161 = _weightQ8_63_12_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_12_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_162 = _weightQ8_63_12_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_12_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_163 = _weightQ8_63_12_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_12_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_164 = _weightQ8_63_12_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_12_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_165 = _weightQ8_63_12_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_12_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_166 = _weightQ8_63_12_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_12_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_167 = _weightQ8_63_12_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_12_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_168 = _weightQ8_63_12_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_12_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_169 = _weightQ8_63_12_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_12_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_170 = _weightQ8_63_12_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_12_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_171 = _weightQ8_63_12_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_12_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_172 = _weightQ8_63_12_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_12_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_173 = _weightQ8_63_12_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_12_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_174 = _weightQ8_63_12_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_12_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_175 = _weightQ8_63_12_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_12_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_176 = _weightQ8_63_12_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_12_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_177 = _weightQ8_63_12_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_12_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_178 = _weightQ8_63_12_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_12_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_179 = _weightQ8_63_12_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_12_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_180 = _weightQ8_63_12_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_12_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_181 = _weightQ8_63_12_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_12_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_182 = _weightQ8_63_12_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_12_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_183 = _weightQ8_63_12_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_12_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_184 = _weightQ8_63_12_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_12_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_185 = _weightQ8_63_12_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_12_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_186 = _weightQ8_63_12_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_12_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_187 = _weightQ8_63_12_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_12_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_188 = _weightQ8_63_12_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_12_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_leadingZeros_T_189 = _weightQ8_63_12_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_12_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_12_leadingZeros = _weightQ8_63_12_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_12_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_12_expRaw_T_1 = 6'h1f - weightQ8_63_12_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_12_expRaw = weightQ8_63_12_isZero ? 6'h0 : _weightQ8_63_12_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_12_shiftAmt_T_2 = weightQ8_63_12_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_12_shiftAmt = weightQ8_63_12_expRaw > 6'h3 ? _weightQ8_63_12_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_12_mantissaRaw_T = weightQ8_63_12_absClipped >> weightQ8_63_12_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_12_mantissaRaw = _weightQ8_63_12_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_12_mantissa = weightQ8_63_12_expRaw >= 6'h3 ? weightQ8_63_12_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_12_expAdjusted = weightQ8_63_12_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_12_exp_T_4 = weightQ8_63_12_expAdjusted > 7'hf ? 4'hf : weightQ8_63_12_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_12_exp = weightQ8_63_12_isZero ? 4'h0 : _weightQ8_63_12_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_12_fp8 = {weightQ8_63_12_clippedX[31],weightQ8_63_12_exp,weightQ8_63_12_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_13_T = {24'h0,linear_weight_63_13}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_13_sign = _weightQ8_63_13_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_13_absX_T = ~_weightQ8_63_13_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_13_absX_T_2 = _weightQ8_63_13_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_13_absX = weightQ8_63_13_sign ? _weightQ8_63_13_absX_T_2 : _weightQ8_63_13_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_13_shiftedX_T_1 = _GEN_14432 - weightQ8_63_13_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_13_shiftedX_T_3 = weightQ8_63_13_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_13_shiftedX = weightQ8_63_13_sign ? _weightQ8_63_13_shiftedX_T_1 :
    _weightQ8_63_13_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_13_scaledX_T_1 = weightQ8_63_13_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_13_scaledX = _weightQ8_63_13_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_13_clippedX_T_2 = weightQ8_63_13_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_13_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_13_clippedX = weightQ8_63_13_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_13_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_13_absClipped_T_1 = ~weightQ8_63_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_13_absClipped_T_3 = _weightQ8_63_13_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_13_absClipped = weightQ8_63_13_clippedX[31] ? _weightQ8_63_13_absClipped_T_3 :
    weightQ8_63_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_13_isZero = weightQ8_63_13_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37457 = {{16'd0}, weightQ8_63_13_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_4 = _GEN_37457 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_6 = {weightQ8_63_13_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_8 = _weightQ8_63_13_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_9 = _weightQ8_63_13_leadingZeros_T_4 | _weightQ8_63_13_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37458 = {{8'd0}, _weightQ8_63_13_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_14 = _GEN_37458 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_16 = {_weightQ8_63_13_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_18 = _weightQ8_63_13_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_19 = _weightQ8_63_13_leadingZeros_T_14 | _weightQ8_63_13_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37459 = {{4'd0}, _weightQ8_63_13_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_24 = _GEN_37459 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_26 = {_weightQ8_63_13_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_28 = _weightQ8_63_13_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_29 = _weightQ8_63_13_leadingZeros_T_24 | _weightQ8_63_13_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37460 = {{2'd0}, _weightQ8_63_13_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_34 = _GEN_37460 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_36 = {_weightQ8_63_13_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_38 = _weightQ8_63_13_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_39 = _weightQ8_63_13_leadingZeros_T_34 | _weightQ8_63_13_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37461 = {{1'd0}, _weightQ8_63_13_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_44 = _GEN_37461 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_46 = {_weightQ8_63_13_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_48 = _weightQ8_63_13_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_13_leadingZeros_T_49 = _weightQ8_63_13_leadingZeros_T_44 | _weightQ8_63_13_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37462 = {{8'd0}, weightQ8_63_13_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_55 = _GEN_37462 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_57 = {weightQ8_63_13_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_59 = _weightQ8_63_13_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_60 = _weightQ8_63_13_leadingZeros_T_55 | _weightQ8_63_13_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37463 = {{4'd0}, _weightQ8_63_13_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_65 = _GEN_37463 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_67 = {_weightQ8_63_13_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_69 = _weightQ8_63_13_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_70 = _weightQ8_63_13_leadingZeros_T_65 | _weightQ8_63_13_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37464 = {{2'd0}, _weightQ8_63_13_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_75 = _GEN_37464 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_77 = {_weightQ8_63_13_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_79 = _weightQ8_63_13_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_80 = _weightQ8_63_13_leadingZeros_T_75 | _weightQ8_63_13_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37465 = {{1'd0}, _weightQ8_63_13_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_85 = _GEN_37465 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_87 = {_weightQ8_63_13_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_89 = _weightQ8_63_13_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_13_leadingZeros_T_90 = _weightQ8_63_13_leadingZeros_T_85 | _weightQ8_63_13_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_13_leadingZeros_T_93 = {_weightQ8_63_13_leadingZeros_T_49,_weightQ8_63_13_leadingZeros_T_90,
    weightQ8_63_13_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_143 = _weightQ8_63_13_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_144 = _weightQ8_63_13_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_13_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_145 = _weightQ8_63_13_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_13_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_146 = _weightQ8_63_13_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_13_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_147 = _weightQ8_63_13_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_13_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_148 = _weightQ8_63_13_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_13_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_149 = _weightQ8_63_13_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_13_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_150 = _weightQ8_63_13_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_13_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_151 = _weightQ8_63_13_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_13_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_152 = _weightQ8_63_13_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_13_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_153 = _weightQ8_63_13_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_13_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_154 = _weightQ8_63_13_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_13_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_155 = _weightQ8_63_13_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_13_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_156 = _weightQ8_63_13_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_13_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_157 = _weightQ8_63_13_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_13_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_158 = _weightQ8_63_13_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_13_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_159 = _weightQ8_63_13_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_13_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_160 = _weightQ8_63_13_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_13_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_161 = _weightQ8_63_13_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_13_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_162 = _weightQ8_63_13_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_13_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_163 = _weightQ8_63_13_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_13_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_164 = _weightQ8_63_13_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_13_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_165 = _weightQ8_63_13_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_13_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_166 = _weightQ8_63_13_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_13_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_167 = _weightQ8_63_13_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_13_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_168 = _weightQ8_63_13_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_13_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_169 = _weightQ8_63_13_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_13_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_170 = _weightQ8_63_13_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_13_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_171 = _weightQ8_63_13_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_13_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_172 = _weightQ8_63_13_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_13_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_173 = _weightQ8_63_13_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_13_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_174 = _weightQ8_63_13_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_13_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_175 = _weightQ8_63_13_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_13_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_176 = _weightQ8_63_13_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_13_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_177 = _weightQ8_63_13_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_13_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_178 = _weightQ8_63_13_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_13_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_179 = _weightQ8_63_13_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_13_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_180 = _weightQ8_63_13_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_13_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_181 = _weightQ8_63_13_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_13_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_182 = _weightQ8_63_13_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_13_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_183 = _weightQ8_63_13_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_13_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_184 = _weightQ8_63_13_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_13_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_185 = _weightQ8_63_13_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_13_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_186 = _weightQ8_63_13_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_13_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_187 = _weightQ8_63_13_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_13_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_188 = _weightQ8_63_13_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_13_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_leadingZeros_T_189 = _weightQ8_63_13_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_13_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_13_leadingZeros = _weightQ8_63_13_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_13_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_13_expRaw_T_1 = 6'h1f - weightQ8_63_13_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_13_expRaw = weightQ8_63_13_isZero ? 6'h0 : _weightQ8_63_13_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_13_shiftAmt_T_2 = weightQ8_63_13_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_13_shiftAmt = weightQ8_63_13_expRaw > 6'h3 ? _weightQ8_63_13_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_13_mantissaRaw_T = weightQ8_63_13_absClipped >> weightQ8_63_13_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_13_mantissaRaw = _weightQ8_63_13_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_13_mantissa = weightQ8_63_13_expRaw >= 6'h3 ? weightQ8_63_13_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_13_expAdjusted = weightQ8_63_13_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_13_exp_T_4 = weightQ8_63_13_expAdjusted > 7'hf ? 4'hf : weightQ8_63_13_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_13_exp = weightQ8_63_13_isZero ? 4'h0 : _weightQ8_63_13_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_13_fp8 = {weightQ8_63_13_clippedX[31],weightQ8_63_13_exp,weightQ8_63_13_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_14_T = {24'h0,linear_weight_63_14}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_14_sign = _weightQ8_63_14_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_14_absX_T = ~_weightQ8_63_14_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_14_absX_T_2 = _weightQ8_63_14_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_14_absX = weightQ8_63_14_sign ? _weightQ8_63_14_absX_T_2 : _weightQ8_63_14_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_14_shiftedX_T_1 = _GEN_14432 - weightQ8_63_14_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_14_shiftedX_T_3 = weightQ8_63_14_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_14_shiftedX = weightQ8_63_14_sign ? _weightQ8_63_14_shiftedX_T_1 :
    _weightQ8_63_14_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_14_scaledX_T_1 = weightQ8_63_14_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_14_scaledX = _weightQ8_63_14_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_14_clippedX_T_2 = weightQ8_63_14_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_14_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_14_clippedX = weightQ8_63_14_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_14_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_14_absClipped_T_1 = ~weightQ8_63_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_14_absClipped_T_3 = _weightQ8_63_14_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_14_absClipped = weightQ8_63_14_clippedX[31] ? _weightQ8_63_14_absClipped_T_3 :
    weightQ8_63_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_14_isZero = weightQ8_63_14_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37468 = {{16'd0}, weightQ8_63_14_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_4 = _GEN_37468 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_6 = {weightQ8_63_14_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_8 = _weightQ8_63_14_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_9 = _weightQ8_63_14_leadingZeros_T_4 | _weightQ8_63_14_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37469 = {{8'd0}, _weightQ8_63_14_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_14 = _GEN_37469 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_16 = {_weightQ8_63_14_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_18 = _weightQ8_63_14_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_19 = _weightQ8_63_14_leadingZeros_T_14 | _weightQ8_63_14_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37470 = {{4'd0}, _weightQ8_63_14_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_24 = _GEN_37470 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_26 = {_weightQ8_63_14_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_28 = _weightQ8_63_14_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_29 = _weightQ8_63_14_leadingZeros_T_24 | _weightQ8_63_14_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37471 = {{2'd0}, _weightQ8_63_14_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_34 = _GEN_37471 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_36 = {_weightQ8_63_14_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_38 = _weightQ8_63_14_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_39 = _weightQ8_63_14_leadingZeros_T_34 | _weightQ8_63_14_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37472 = {{1'd0}, _weightQ8_63_14_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_44 = _GEN_37472 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_46 = {_weightQ8_63_14_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_48 = _weightQ8_63_14_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_14_leadingZeros_T_49 = _weightQ8_63_14_leadingZeros_T_44 | _weightQ8_63_14_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37473 = {{8'd0}, weightQ8_63_14_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_55 = _GEN_37473 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_57 = {weightQ8_63_14_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_59 = _weightQ8_63_14_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_60 = _weightQ8_63_14_leadingZeros_T_55 | _weightQ8_63_14_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37474 = {{4'd0}, _weightQ8_63_14_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_65 = _GEN_37474 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_67 = {_weightQ8_63_14_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_69 = _weightQ8_63_14_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_70 = _weightQ8_63_14_leadingZeros_T_65 | _weightQ8_63_14_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37475 = {{2'd0}, _weightQ8_63_14_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_75 = _GEN_37475 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_77 = {_weightQ8_63_14_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_79 = _weightQ8_63_14_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_80 = _weightQ8_63_14_leadingZeros_T_75 | _weightQ8_63_14_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37476 = {{1'd0}, _weightQ8_63_14_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_85 = _GEN_37476 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_87 = {_weightQ8_63_14_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_89 = _weightQ8_63_14_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_14_leadingZeros_T_90 = _weightQ8_63_14_leadingZeros_T_85 | _weightQ8_63_14_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_14_leadingZeros_T_93 = {_weightQ8_63_14_leadingZeros_T_49,_weightQ8_63_14_leadingZeros_T_90,
    weightQ8_63_14_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_143 = _weightQ8_63_14_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_144 = _weightQ8_63_14_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_14_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_145 = _weightQ8_63_14_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_14_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_146 = _weightQ8_63_14_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_14_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_147 = _weightQ8_63_14_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_14_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_148 = _weightQ8_63_14_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_14_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_149 = _weightQ8_63_14_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_14_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_150 = _weightQ8_63_14_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_14_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_151 = _weightQ8_63_14_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_14_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_152 = _weightQ8_63_14_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_14_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_153 = _weightQ8_63_14_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_14_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_154 = _weightQ8_63_14_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_14_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_155 = _weightQ8_63_14_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_14_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_156 = _weightQ8_63_14_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_14_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_157 = _weightQ8_63_14_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_14_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_158 = _weightQ8_63_14_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_14_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_159 = _weightQ8_63_14_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_14_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_160 = _weightQ8_63_14_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_14_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_161 = _weightQ8_63_14_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_14_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_162 = _weightQ8_63_14_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_14_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_163 = _weightQ8_63_14_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_14_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_164 = _weightQ8_63_14_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_14_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_165 = _weightQ8_63_14_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_14_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_166 = _weightQ8_63_14_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_14_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_167 = _weightQ8_63_14_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_14_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_168 = _weightQ8_63_14_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_14_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_169 = _weightQ8_63_14_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_14_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_170 = _weightQ8_63_14_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_14_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_171 = _weightQ8_63_14_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_14_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_172 = _weightQ8_63_14_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_14_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_173 = _weightQ8_63_14_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_14_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_174 = _weightQ8_63_14_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_14_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_175 = _weightQ8_63_14_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_14_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_176 = _weightQ8_63_14_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_14_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_177 = _weightQ8_63_14_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_14_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_178 = _weightQ8_63_14_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_14_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_179 = _weightQ8_63_14_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_14_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_180 = _weightQ8_63_14_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_14_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_181 = _weightQ8_63_14_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_14_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_182 = _weightQ8_63_14_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_14_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_183 = _weightQ8_63_14_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_14_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_184 = _weightQ8_63_14_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_14_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_185 = _weightQ8_63_14_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_14_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_186 = _weightQ8_63_14_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_14_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_187 = _weightQ8_63_14_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_14_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_188 = _weightQ8_63_14_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_14_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_leadingZeros_T_189 = _weightQ8_63_14_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_14_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_14_leadingZeros = _weightQ8_63_14_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_14_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_14_expRaw_T_1 = 6'h1f - weightQ8_63_14_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_14_expRaw = weightQ8_63_14_isZero ? 6'h0 : _weightQ8_63_14_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_14_shiftAmt_T_2 = weightQ8_63_14_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_14_shiftAmt = weightQ8_63_14_expRaw > 6'h3 ? _weightQ8_63_14_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_14_mantissaRaw_T = weightQ8_63_14_absClipped >> weightQ8_63_14_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_14_mantissaRaw = _weightQ8_63_14_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_14_mantissa = weightQ8_63_14_expRaw >= 6'h3 ? weightQ8_63_14_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_14_expAdjusted = weightQ8_63_14_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_14_exp_T_4 = weightQ8_63_14_expAdjusted > 7'hf ? 4'hf : weightQ8_63_14_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_14_exp = weightQ8_63_14_isZero ? 4'h0 : _weightQ8_63_14_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_14_fp8 = {weightQ8_63_14_clippedX[31],weightQ8_63_14_exp,weightQ8_63_14_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_15_T = {24'h0,linear_weight_63_15}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_15_sign = _weightQ8_63_15_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_15_absX_T = ~_weightQ8_63_15_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_15_absX_T_2 = _weightQ8_63_15_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_15_absX = weightQ8_63_15_sign ? _weightQ8_63_15_absX_T_2 : _weightQ8_63_15_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_15_shiftedX_T_1 = _GEN_14432 - weightQ8_63_15_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_15_shiftedX_T_3 = weightQ8_63_15_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_15_shiftedX = weightQ8_63_15_sign ? _weightQ8_63_15_shiftedX_T_1 :
    _weightQ8_63_15_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_15_scaledX_T_1 = weightQ8_63_15_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_15_scaledX = _weightQ8_63_15_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_15_clippedX_T_2 = weightQ8_63_15_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_15_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_15_clippedX = weightQ8_63_15_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_15_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_15_absClipped_T_1 = ~weightQ8_63_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_15_absClipped_T_3 = _weightQ8_63_15_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_15_absClipped = weightQ8_63_15_clippedX[31] ? _weightQ8_63_15_absClipped_T_3 :
    weightQ8_63_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_15_isZero = weightQ8_63_15_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37479 = {{16'd0}, weightQ8_63_15_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_4 = _GEN_37479 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_6 = {weightQ8_63_15_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_8 = _weightQ8_63_15_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_9 = _weightQ8_63_15_leadingZeros_T_4 | _weightQ8_63_15_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37480 = {{8'd0}, _weightQ8_63_15_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_14 = _GEN_37480 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_16 = {_weightQ8_63_15_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_18 = _weightQ8_63_15_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_19 = _weightQ8_63_15_leadingZeros_T_14 | _weightQ8_63_15_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37481 = {{4'd0}, _weightQ8_63_15_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_24 = _GEN_37481 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_26 = {_weightQ8_63_15_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_28 = _weightQ8_63_15_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_29 = _weightQ8_63_15_leadingZeros_T_24 | _weightQ8_63_15_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37482 = {{2'd0}, _weightQ8_63_15_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_34 = _GEN_37482 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_36 = {_weightQ8_63_15_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_38 = _weightQ8_63_15_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_39 = _weightQ8_63_15_leadingZeros_T_34 | _weightQ8_63_15_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37483 = {{1'd0}, _weightQ8_63_15_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_44 = _GEN_37483 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_46 = {_weightQ8_63_15_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_48 = _weightQ8_63_15_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_15_leadingZeros_T_49 = _weightQ8_63_15_leadingZeros_T_44 | _weightQ8_63_15_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37484 = {{8'd0}, weightQ8_63_15_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_55 = _GEN_37484 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_57 = {weightQ8_63_15_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_59 = _weightQ8_63_15_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_60 = _weightQ8_63_15_leadingZeros_T_55 | _weightQ8_63_15_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37485 = {{4'd0}, _weightQ8_63_15_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_65 = _GEN_37485 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_67 = {_weightQ8_63_15_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_69 = _weightQ8_63_15_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_70 = _weightQ8_63_15_leadingZeros_T_65 | _weightQ8_63_15_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37486 = {{2'd0}, _weightQ8_63_15_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_75 = _GEN_37486 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_77 = {_weightQ8_63_15_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_79 = _weightQ8_63_15_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_80 = _weightQ8_63_15_leadingZeros_T_75 | _weightQ8_63_15_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37487 = {{1'd0}, _weightQ8_63_15_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_85 = _GEN_37487 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_87 = {_weightQ8_63_15_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_89 = _weightQ8_63_15_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_15_leadingZeros_T_90 = _weightQ8_63_15_leadingZeros_T_85 | _weightQ8_63_15_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_15_leadingZeros_T_93 = {_weightQ8_63_15_leadingZeros_T_49,_weightQ8_63_15_leadingZeros_T_90,
    weightQ8_63_15_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_143 = _weightQ8_63_15_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_144 = _weightQ8_63_15_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_15_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_145 = _weightQ8_63_15_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_15_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_146 = _weightQ8_63_15_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_15_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_147 = _weightQ8_63_15_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_15_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_148 = _weightQ8_63_15_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_15_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_149 = _weightQ8_63_15_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_15_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_150 = _weightQ8_63_15_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_15_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_151 = _weightQ8_63_15_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_15_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_152 = _weightQ8_63_15_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_15_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_153 = _weightQ8_63_15_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_15_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_154 = _weightQ8_63_15_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_15_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_155 = _weightQ8_63_15_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_15_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_156 = _weightQ8_63_15_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_15_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_157 = _weightQ8_63_15_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_15_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_158 = _weightQ8_63_15_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_15_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_159 = _weightQ8_63_15_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_15_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_160 = _weightQ8_63_15_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_15_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_161 = _weightQ8_63_15_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_15_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_162 = _weightQ8_63_15_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_15_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_163 = _weightQ8_63_15_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_15_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_164 = _weightQ8_63_15_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_15_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_165 = _weightQ8_63_15_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_15_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_166 = _weightQ8_63_15_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_15_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_167 = _weightQ8_63_15_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_15_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_168 = _weightQ8_63_15_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_15_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_169 = _weightQ8_63_15_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_15_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_170 = _weightQ8_63_15_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_15_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_171 = _weightQ8_63_15_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_15_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_172 = _weightQ8_63_15_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_15_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_173 = _weightQ8_63_15_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_15_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_174 = _weightQ8_63_15_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_15_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_175 = _weightQ8_63_15_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_15_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_176 = _weightQ8_63_15_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_15_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_177 = _weightQ8_63_15_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_15_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_178 = _weightQ8_63_15_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_15_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_179 = _weightQ8_63_15_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_15_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_180 = _weightQ8_63_15_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_15_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_181 = _weightQ8_63_15_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_15_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_182 = _weightQ8_63_15_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_15_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_183 = _weightQ8_63_15_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_15_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_184 = _weightQ8_63_15_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_15_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_185 = _weightQ8_63_15_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_15_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_186 = _weightQ8_63_15_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_15_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_187 = _weightQ8_63_15_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_15_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_188 = _weightQ8_63_15_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_15_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_leadingZeros_T_189 = _weightQ8_63_15_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_15_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_15_leadingZeros = _weightQ8_63_15_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_15_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_15_expRaw_T_1 = 6'h1f - weightQ8_63_15_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_15_expRaw = weightQ8_63_15_isZero ? 6'h0 : _weightQ8_63_15_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_15_shiftAmt_T_2 = weightQ8_63_15_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_15_shiftAmt = weightQ8_63_15_expRaw > 6'h3 ? _weightQ8_63_15_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_15_mantissaRaw_T = weightQ8_63_15_absClipped >> weightQ8_63_15_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_15_mantissaRaw = _weightQ8_63_15_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_15_mantissa = weightQ8_63_15_expRaw >= 6'h3 ? weightQ8_63_15_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_15_expAdjusted = weightQ8_63_15_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_15_exp_T_4 = weightQ8_63_15_expAdjusted > 7'hf ? 4'hf : weightQ8_63_15_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_15_exp = weightQ8_63_15_isZero ? 4'h0 : _weightQ8_63_15_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_15_fp8 = {weightQ8_63_15_clippedX[31],weightQ8_63_15_exp,weightQ8_63_15_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_16_T = {24'h0,linear_weight_63_16}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_16_sign = _weightQ8_63_16_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_16_absX_T = ~_weightQ8_63_16_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_16_absX_T_2 = _weightQ8_63_16_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_16_absX = weightQ8_63_16_sign ? _weightQ8_63_16_absX_T_2 : _weightQ8_63_16_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_16_shiftedX_T_1 = _GEN_14432 - weightQ8_63_16_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_16_shiftedX_T_3 = weightQ8_63_16_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_16_shiftedX = weightQ8_63_16_sign ? _weightQ8_63_16_shiftedX_T_1 :
    _weightQ8_63_16_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_16_scaledX_T_1 = weightQ8_63_16_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_16_scaledX = _weightQ8_63_16_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_16_clippedX_T_2 = weightQ8_63_16_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_16_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_16_clippedX = weightQ8_63_16_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_16_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_16_absClipped_T_1 = ~weightQ8_63_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_16_absClipped_T_3 = _weightQ8_63_16_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_16_absClipped = weightQ8_63_16_clippedX[31] ? _weightQ8_63_16_absClipped_T_3 :
    weightQ8_63_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_16_isZero = weightQ8_63_16_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37490 = {{16'd0}, weightQ8_63_16_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_4 = _GEN_37490 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_6 = {weightQ8_63_16_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_8 = _weightQ8_63_16_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_9 = _weightQ8_63_16_leadingZeros_T_4 | _weightQ8_63_16_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37491 = {{8'd0}, _weightQ8_63_16_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_14 = _GEN_37491 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_16 = {_weightQ8_63_16_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_18 = _weightQ8_63_16_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_19 = _weightQ8_63_16_leadingZeros_T_14 | _weightQ8_63_16_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37492 = {{4'd0}, _weightQ8_63_16_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_24 = _GEN_37492 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_26 = {_weightQ8_63_16_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_28 = _weightQ8_63_16_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_29 = _weightQ8_63_16_leadingZeros_T_24 | _weightQ8_63_16_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37493 = {{2'd0}, _weightQ8_63_16_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_34 = _GEN_37493 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_36 = {_weightQ8_63_16_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_38 = _weightQ8_63_16_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_39 = _weightQ8_63_16_leadingZeros_T_34 | _weightQ8_63_16_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37494 = {{1'd0}, _weightQ8_63_16_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_44 = _GEN_37494 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_46 = {_weightQ8_63_16_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_48 = _weightQ8_63_16_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_16_leadingZeros_T_49 = _weightQ8_63_16_leadingZeros_T_44 | _weightQ8_63_16_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37495 = {{8'd0}, weightQ8_63_16_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_55 = _GEN_37495 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_57 = {weightQ8_63_16_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_59 = _weightQ8_63_16_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_60 = _weightQ8_63_16_leadingZeros_T_55 | _weightQ8_63_16_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37496 = {{4'd0}, _weightQ8_63_16_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_65 = _GEN_37496 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_67 = {_weightQ8_63_16_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_69 = _weightQ8_63_16_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_70 = _weightQ8_63_16_leadingZeros_T_65 | _weightQ8_63_16_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37497 = {{2'd0}, _weightQ8_63_16_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_75 = _GEN_37497 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_77 = {_weightQ8_63_16_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_79 = _weightQ8_63_16_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_80 = _weightQ8_63_16_leadingZeros_T_75 | _weightQ8_63_16_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37498 = {{1'd0}, _weightQ8_63_16_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_85 = _GEN_37498 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_87 = {_weightQ8_63_16_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_89 = _weightQ8_63_16_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_16_leadingZeros_T_90 = _weightQ8_63_16_leadingZeros_T_85 | _weightQ8_63_16_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_16_leadingZeros_T_93 = {_weightQ8_63_16_leadingZeros_T_49,_weightQ8_63_16_leadingZeros_T_90,
    weightQ8_63_16_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_143 = _weightQ8_63_16_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_144 = _weightQ8_63_16_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_16_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_145 = _weightQ8_63_16_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_16_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_146 = _weightQ8_63_16_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_16_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_147 = _weightQ8_63_16_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_16_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_148 = _weightQ8_63_16_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_16_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_149 = _weightQ8_63_16_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_16_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_150 = _weightQ8_63_16_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_16_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_151 = _weightQ8_63_16_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_16_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_152 = _weightQ8_63_16_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_16_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_153 = _weightQ8_63_16_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_16_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_154 = _weightQ8_63_16_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_16_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_155 = _weightQ8_63_16_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_16_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_156 = _weightQ8_63_16_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_16_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_157 = _weightQ8_63_16_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_16_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_158 = _weightQ8_63_16_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_16_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_159 = _weightQ8_63_16_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_16_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_160 = _weightQ8_63_16_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_16_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_161 = _weightQ8_63_16_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_16_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_162 = _weightQ8_63_16_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_16_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_163 = _weightQ8_63_16_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_16_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_164 = _weightQ8_63_16_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_16_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_165 = _weightQ8_63_16_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_16_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_166 = _weightQ8_63_16_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_16_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_167 = _weightQ8_63_16_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_16_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_168 = _weightQ8_63_16_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_16_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_169 = _weightQ8_63_16_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_16_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_170 = _weightQ8_63_16_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_16_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_171 = _weightQ8_63_16_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_16_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_172 = _weightQ8_63_16_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_16_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_173 = _weightQ8_63_16_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_16_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_174 = _weightQ8_63_16_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_16_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_175 = _weightQ8_63_16_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_16_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_176 = _weightQ8_63_16_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_16_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_177 = _weightQ8_63_16_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_16_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_178 = _weightQ8_63_16_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_16_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_179 = _weightQ8_63_16_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_16_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_180 = _weightQ8_63_16_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_16_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_181 = _weightQ8_63_16_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_16_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_182 = _weightQ8_63_16_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_16_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_183 = _weightQ8_63_16_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_16_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_184 = _weightQ8_63_16_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_16_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_185 = _weightQ8_63_16_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_16_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_186 = _weightQ8_63_16_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_16_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_187 = _weightQ8_63_16_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_16_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_188 = _weightQ8_63_16_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_16_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_leadingZeros_T_189 = _weightQ8_63_16_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_16_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_16_leadingZeros = _weightQ8_63_16_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_16_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_16_expRaw_T_1 = 6'h1f - weightQ8_63_16_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_16_expRaw = weightQ8_63_16_isZero ? 6'h0 : _weightQ8_63_16_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_16_shiftAmt_T_2 = weightQ8_63_16_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_16_shiftAmt = weightQ8_63_16_expRaw > 6'h3 ? _weightQ8_63_16_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_16_mantissaRaw_T = weightQ8_63_16_absClipped >> weightQ8_63_16_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_16_mantissaRaw = _weightQ8_63_16_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_16_mantissa = weightQ8_63_16_expRaw >= 6'h3 ? weightQ8_63_16_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_16_expAdjusted = weightQ8_63_16_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_16_exp_T_4 = weightQ8_63_16_expAdjusted > 7'hf ? 4'hf : weightQ8_63_16_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_16_exp = weightQ8_63_16_isZero ? 4'h0 : _weightQ8_63_16_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_16_fp8 = {weightQ8_63_16_clippedX[31],weightQ8_63_16_exp,weightQ8_63_16_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_17_T = {24'h0,linear_weight_63_17}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_17_sign = _weightQ8_63_17_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_17_absX_T = ~_weightQ8_63_17_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_17_absX_T_2 = _weightQ8_63_17_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_17_absX = weightQ8_63_17_sign ? _weightQ8_63_17_absX_T_2 : _weightQ8_63_17_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_17_shiftedX_T_1 = _GEN_14432 - weightQ8_63_17_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_17_shiftedX_T_3 = weightQ8_63_17_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_17_shiftedX = weightQ8_63_17_sign ? _weightQ8_63_17_shiftedX_T_1 :
    _weightQ8_63_17_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_17_scaledX_T_1 = weightQ8_63_17_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_17_scaledX = _weightQ8_63_17_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_17_clippedX_T_2 = weightQ8_63_17_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_17_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_17_clippedX = weightQ8_63_17_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_17_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_17_absClipped_T_1 = ~weightQ8_63_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_17_absClipped_T_3 = _weightQ8_63_17_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_17_absClipped = weightQ8_63_17_clippedX[31] ? _weightQ8_63_17_absClipped_T_3 :
    weightQ8_63_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_17_isZero = weightQ8_63_17_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37501 = {{16'd0}, weightQ8_63_17_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_4 = _GEN_37501 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_6 = {weightQ8_63_17_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_8 = _weightQ8_63_17_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_9 = _weightQ8_63_17_leadingZeros_T_4 | _weightQ8_63_17_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37502 = {{8'd0}, _weightQ8_63_17_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_14 = _GEN_37502 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_16 = {_weightQ8_63_17_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_18 = _weightQ8_63_17_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_19 = _weightQ8_63_17_leadingZeros_T_14 | _weightQ8_63_17_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37503 = {{4'd0}, _weightQ8_63_17_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_24 = _GEN_37503 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_26 = {_weightQ8_63_17_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_28 = _weightQ8_63_17_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_29 = _weightQ8_63_17_leadingZeros_T_24 | _weightQ8_63_17_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37504 = {{2'd0}, _weightQ8_63_17_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_34 = _GEN_37504 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_36 = {_weightQ8_63_17_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_38 = _weightQ8_63_17_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_39 = _weightQ8_63_17_leadingZeros_T_34 | _weightQ8_63_17_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37505 = {{1'd0}, _weightQ8_63_17_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_44 = _GEN_37505 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_46 = {_weightQ8_63_17_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_48 = _weightQ8_63_17_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_17_leadingZeros_T_49 = _weightQ8_63_17_leadingZeros_T_44 | _weightQ8_63_17_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37506 = {{8'd0}, weightQ8_63_17_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_55 = _GEN_37506 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_57 = {weightQ8_63_17_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_59 = _weightQ8_63_17_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_60 = _weightQ8_63_17_leadingZeros_T_55 | _weightQ8_63_17_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37507 = {{4'd0}, _weightQ8_63_17_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_65 = _GEN_37507 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_67 = {_weightQ8_63_17_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_69 = _weightQ8_63_17_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_70 = _weightQ8_63_17_leadingZeros_T_65 | _weightQ8_63_17_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37508 = {{2'd0}, _weightQ8_63_17_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_75 = _GEN_37508 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_77 = {_weightQ8_63_17_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_79 = _weightQ8_63_17_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_80 = _weightQ8_63_17_leadingZeros_T_75 | _weightQ8_63_17_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37509 = {{1'd0}, _weightQ8_63_17_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_85 = _GEN_37509 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_87 = {_weightQ8_63_17_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_89 = _weightQ8_63_17_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_17_leadingZeros_T_90 = _weightQ8_63_17_leadingZeros_T_85 | _weightQ8_63_17_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_17_leadingZeros_T_93 = {_weightQ8_63_17_leadingZeros_T_49,_weightQ8_63_17_leadingZeros_T_90,
    weightQ8_63_17_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_143 = _weightQ8_63_17_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_144 = _weightQ8_63_17_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_17_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_145 = _weightQ8_63_17_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_17_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_146 = _weightQ8_63_17_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_17_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_147 = _weightQ8_63_17_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_17_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_148 = _weightQ8_63_17_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_17_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_149 = _weightQ8_63_17_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_17_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_150 = _weightQ8_63_17_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_17_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_151 = _weightQ8_63_17_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_17_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_152 = _weightQ8_63_17_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_17_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_153 = _weightQ8_63_17_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_17_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_154 = _weightQ8_63_17_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_17_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_155 = _weightQ8_63_17_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_17_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_156 = _weightQ8_63_17_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_17_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_157 = _weightQ8_63_17_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_17_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_158 = _weightQ8_63_17_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_17_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_159 = _weightQ8_63_17_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_17_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_160 = _weightQ8_63_17_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_17_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_161 = _weightQ8_63_17_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_17_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_162 = _weightQ8_63_17_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_17_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_163 = _weightQ8_63_17_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_17_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_164 = _weightQ8_63_17_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_17_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_165 = _weightQ8_63_17_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_17_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_166 = _weightQ8_63_17_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_17_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_167 = _weightQ8_63_17_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_17_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_168 = _weightQ8_63_17_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_17_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_169 = _weightQ8_63_17_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_17_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_170 = _weightQ8_63_17_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_17_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_171 = _weightQ8_63_17_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_17_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_172 = _weightQ8_63_17_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_17_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_173 = _weightQ8_63_17_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_17_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_174 = _weightQ8_63_17_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_17_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_175 = _weightQ8_63_17_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_17_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_176 = _weightQ8_63_17_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_17_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_177 = _weightQ8_63_17_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_17_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_178 = _weightQ8_63_17_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_17_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_179 = _weightQ8_63_17_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_17_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_180 = _weightQ8_63_17_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_17_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_181 = _weightQ8_63_17_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_17_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_182 = _weightQ8_63_17_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_17_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_183 = _weightQ8_63_17_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_17_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_184 = _weightQ8_63_17_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_17_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_185 = _weightQ8_63_17_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_17_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_186 = _weightQ8_63_17_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_17_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_187 = _weightQ8_63_17_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_17_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_188 = _weightQ8_63_17_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_17_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_leadingZeros_T_189 = _weightQ8_63_17_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_17_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_17_leadingZeros = _weightQ8_63_17_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_17_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_17_expRaw_T_1 = 6'h1f - weightQ8_63_17_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_17_expRaw = weightQ8_63_17_isZero ? 6'h0 : _weightQ8_63_17_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_17_shiftAmt_T_2 = weightQ8_63_17_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_17_shiftAmt = weightQ8_63_17_expRaw > 6'h3 ? _weightQ8_63_17_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_17_mantissaRaw_T = weightQ8_63_17_absClipped >> weightQ8_63_17_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_17_mantissaRaw = _weightQ8_63_17_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_17_mantissa = weightQ8_63_17_expRaw >= 6'h3 ? weightQ8_63_17_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_17_expAdjusted = weightQ8_63_17_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_17_exp_T_4 = weightQ8_63_17_expAdjusted > 7'hf ? 4'hf : weightQ8_63_17_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_17_exp = weightQ8_63_17_isZero ? 4'h0 : _weightQ8_63_17_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_17_fp8 = {weightQ8_63_17_clippedX[31],weightQ8_63_17_exp,weightQ8_63_17_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_18_T = {24'h0,linear_weight_63_18}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_18_sign = _weightQ8_63_18_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_18_absX_T = ~_weightQ8_63_18_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_18_absX_T_2 = _weightQ8_63_18_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_18_absX = weightQ8_63_18_sign ? _weightQ8_63_18_absX_T_2 : _weightQ8_63_18_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_18_shiftedX_T_1 = _GEN_14432 - weightQ8_63_18_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_18_shiftedX_T_3 = weightQ8_63_18_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_18_shiftedX = weightQ8_63_18_sign ? _weightQ8_63_18_shiftedX_T_1 :
    _weightQ8_63_18_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_18_scaledX_T_1 = weightQ8_63_18_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_18_scaledX = _weightQ8_63_18_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_18_clippedX_T_2 = weightQ8_63_18_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_18_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_18_clippedX = weightQ8_63_18_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_18_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_18_absClipped_T_1 = ~weightQ8_63_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_18_absClipped_T_3 = _weightQ8_63_18_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_18_absClipped = weightQ8_63_18_clippedX[31] ? _weightQ8_63_18_absClipped_T_3 :
    weightQ8_63_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_18_isZero = weightQ8_63_18_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37512 = {{16'd0}, weightQ8_63_18_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_4 = _GEN_37512 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_6 = {weightQ8_63_18_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_8 = _weightQ8_63_18_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_9 = _weightQ8_63_18_leadingZeros_T_4 | _weightQ8_63_18_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37513 = {{8'd0}, _weightQ8_63_18_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_14 = _GEN_37513 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_16 = {_weightQ8_63_18_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_18 = _weightQ8_63_18_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_19 = _weightQ8_63_18_leadingZeros_T_14 | _weightQ8_63_18_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37514 = {{4'd0}, _weightQ8_63_18_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_24 = _GEN_37514 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_26 = {_weightQ8_63_18_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_28 = _weightQ8_63_18_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_29 = _weightQ8_63_18_leadingZeros_T_24 | _weightQ8_63_18_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37515 = {{2'd0}, _weightQ8_63_18_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_34 = _GEN_37515 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_36 = {_weightQ8_63_18_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_38 = _weightQ8_63_18_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_39 = _weightQ8_63_18_leadingZeros_T_34 | _weightQ8_63_18_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37516 = {{1'd0}, _weightQ8_63_18_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_44 = _GEN_37516 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_46 = {_weightQ8_63_18_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_48 = _weightQ8_63_18_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_18_leadingZeros_T_49 = _weightQ8_63_18_leadingZeros_T_44 | _weightQ8_63_18_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37517 = {{8'd0}, weightQ8_63_18_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_55 = _GEN_37517 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_57 = {weightQ8_63_18_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_59 = _weightQ8_63_18_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_60 = _weightQ8_63_18_leadingZeros_T_55 | _weightQ8_63_18_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37518 = {{4'd0}, _weightQ8_63_18_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_65 = _GEN_37518 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_67 = {_weightQ8_63_18_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_69 = _weightQ8_63_18_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_70 = _weightQ8_63_18_leadingZeros_T_65 | _weightQ8_63_18_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37519 = {{2'd0}, _weightQ8_63_18_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_75 = _GEN_37519 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_77 = {_weightQ8_63_18_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_79 = _weightQ8_63_18_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_80 = _weightQ8_63_18_leadingZeros_T_75 | _weightQ8_63_18_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37520 = {{1'd0}, _weightQ8_63_18_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_85 = _GEN_37520 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_87 = {_weightQ8_63_18_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_89 = _weightQ8_63_18_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_18_leadingZeros_T_90 = _weightQ8_63_18_leadingZeros_T_85 | _weightQ8_63_18_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_18_leadingZeros_T_93 = {_weightQ8_63_18_leadingZeros_T_49,_weightQ8_63_18_leadingZeros_T_90,
    weightQ8_63_18_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_143 = _weightQ8_63_18_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_144 = _weightQ8_63_18_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_18_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_145 = _weightQ8_63_18_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_18_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_146 = _weightQ8_63_18_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_18_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_147 = _weightQ8_63_18_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_18_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_148 = _weightQ8_63_18_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_18_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_149 = _weightQ8_63_18_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_18_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_150 = _weightQ8_63_18_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_18_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_151 = _weightQ8_63_18_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_18_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_152 = _weightQ8_63_18_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_18_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_153 = _weightQ8_63_18_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_18_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_154 = _weightQ8_63_18_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_18_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_155 = _weightQ8_63_18_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_18_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_156 = _weightQ8_63_18_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_18_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_157 = _weightQ8_63_18_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_18_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_158 = _weightQ8_63_18_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_18_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_159 = _weightQ8_63_18_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_18_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_160 = _weightQ8_63_18_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_18_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_161 = _weightQ8_63_18_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_18_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_162 = _weightQ8_63_18_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_18_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_163 = _weightQ8_63_18_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_18_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_164 = _weightQ8_63_18_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_18_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_165 = _weightQ8_63_18_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_18_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_166 = _weightQ8_63_18_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_18_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_167 = _weightQ8_63_18_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_18_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_168 = _weightQ8_63_18_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_18_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_169 = _weightQ8_63_18_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_18_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_170 = _weightQ8_63_18_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_18_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_171 = _weightQ8_63_18_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_18_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_172 = _weightQ8_63_18_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_18_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_173 = _weightQ8_63_18_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_18_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_174 = _weightQ8_63_18_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_18_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_175 = _weightQ8_63_18_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_18_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_176 = _weightQ8_63_18_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_18_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_177 = _weightQ8_63_18_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_18_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_178 = _weightQ8_63_18_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_18_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_179 = _weightQ8_63_18_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_18_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_180 = _weightQ8_63_18_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_18_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_181 = _weightQ8_63_18_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_18_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_182 = _weightQ8_63_18_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_18_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_183 = _weightQ8_63_18_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_18_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_184 = _weightQ8_63_18_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_18_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_185 = _weightQ8_63_18_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_18_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_186 = _weightQ8_63_18_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_18_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_187 = _weightQ8_63_18_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_18_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_188 = _weightQ8_63_18_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_18_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_leadingZeros_T_189 = _weightQ8_63_18_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_18_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_18_leadingZeros = _weightQ8_63_18_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_18_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_18_expRaw_T_1 = 6'h1f - weightQ8_63_18_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_18_expRaw = weightQ8_63_18_isZero ? 6'h0 : _weightQ8_63_18_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_18_shiftAmt_T_2 = weightQ8_63_18_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_18_shiftAmt = weightQ8_63_18_expRaw > 6'h3 ? _weightQ8_63_18_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_18_mantissaRaw_T = weightQ8_63_18_absClipped >> weightQ8_63_18_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_18_mantissaRaw = _weightQ8_63_18_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_18_mantissa = weightQ8_63_18_expRaw >= 6'h3 ? weightQ8_63_18_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_18_expAdjusted = weightQ8_63_18_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_18_exp_T_4 = weightQ8_63_18_expAdjusted > 7'hf ? 4'hf : weightQ8_63_18_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_18_exp = weightQ8_63_18_isZero ? 4'h0 : _weightQ8_63_18_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_18_fp8 = {weightQ8_63_18_clippedX[31],weightQ8_63_18_exp,weightQ8_63_18_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_19_T = {24'h0,linear_weight_63_19}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_19_sign = _weightQ8_63_19_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_19_absX_T = ~_weightQ8_63_19_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_19_absX_T_2 = _weightQ8_63_19_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_19_absX = weightQ8_63_19_sign ? _weightQ8_63_19_absX_T_2 : _weightQ8_63_19_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_19_shiftedX_T_1 = _GEN_14432 - weightQ8_63_19_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_19_shiftedX_T_3 = weightQ8_63_19_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_19_shiftedX = weightQ8_63_19_sign ? _weightQ8_63_19_shiftedX_T_1 :
    _weightQ8_63_19_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_19_scaledX_T_1 = weightQ8_63_19_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_19_scaledX = _weightQ8_63_19_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_19_clippedX_T_2 = weightQ8_63_19_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_19_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_19_clippedX = weightQ8_63_19_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_19_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_19_absClipped_T_1 = ~weightQ8_63_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_19_absClipped_T_3 = _weightQ8_63_19_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_19_absClipped = weightQ8_63_19_clippedX[31] ? _weightQ8_63_19_absClipped_T_3 :
    weightQ8_63_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_19_isZero = weightQ8_63_19_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37523 = {{16'd0}, weightQ8_63_19_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_4 = _GEN_37523 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_6 = {weightQ8_63_19_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_8 = _weightQ8_63_19_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_9 = _weightQ8_63_19_leadingZeros_T_4 | _weightQ8_63_19_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37524 = {{8'd0}, _weightQ8_63_19_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_14 = _GEN_37524 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_16 = {_weightQ8_63_19_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_18 = _weightQ8_63_19_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_19 = _weightQ8_63_19_leadingZeros_T_14 | _weightQ8_63_19_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37525 = {{4'd0}, _weightQ8_63_19_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_24 = _GEN_37525 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_26 = {_weightQ8_63_19_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_28 = _weightQ8_63_19_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_29 = _weightQ8_63_19_leadingZeros_T_24 | _weightQ8_63_19_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37526 = {{2'd0}, _weightQ8_63_19_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_34 = _GEN_37526 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_36 = {_weightQ8_63_19_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_38 = _weightQ8_63_19_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_39 = _weightQ8_63_19_leadingZeros_T_34 | _weightQ8_63_19_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37527 = {{1'd0}, _weightQ8_63_19_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_44 = _GEN_37527 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_46 = {_weightQ8_63_19_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_48 = _weightQ8_63_19_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_19_leadingZeros_T_49 = _weightQ8_63_19_leadingZeros_T_44 | _weightQ8_63_19_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37528 = {{8'd0}, weightQ8_63_19_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_55 = _GEN_37528 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_57 = {weightQ8_63_19_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_59 = _weightQ8_63_19_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_60 = _weightQ8_63_19_leadingZeros_T_55 | _weightQ8_63_19_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37529 = {{4'd0}, _weightQ8_63_19_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_65 = _GEN_37529 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_67 = {_weightQ8_63_19_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_69 = _weightQ8_63_19_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_70 = _weightQ8_63_19_leadingZeros_T_65 | _weightQ8_63_19_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37530 = {{2'd0}, _weightQ8_63_19_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_75 = _GEN_37530 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_77 = {_weightQ8_63_19_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_79 = _weightQ8_63_19_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_80 = _weightQ8_63_19_leadingZeros_T_75 | _weightQ8_63_19_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37531 = {{1'd0}, _weightQ8_63_19_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_85 = _GEN_37531 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_87 = {_weightQ8_63_19_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_89 = _weightQ8_63_19_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_19_leadingZeros_T_90 = _weightQ8_63_19_leadingZeros_T_85 | _weightQ8_63_19_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_19_leadingZeros_T_93 = {_weightQ8_63_19_leadingZeros_T_49,_weightQ8_63_19_leadingZeros_T_90,
    weightQ8_63_19_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_143 = _weightQ8_63_19_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_144 = _weightQ8_63_19_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_19_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_145 = _weightQ8_63_19_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_19_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_146 = _weightQ8_63_19_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_19_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_147 = _weightQ8_63_19_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_19_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_148 = _weightQ8_63_19_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_19_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_149 = _weightQ8_63_19_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_19_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_150 = _weightQ8_63_19_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_19_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_151 = _weightQ8_63_19_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_19_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_152 = _weightQ8_63_19_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_19_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_153 = _weightQ8_63_19_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_19_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_154 = _weightQ8_63_19_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_19_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_155 = _weightQ8_63_19_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_19_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_156 = _weightQ8_63_19_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_19_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_157 = _weightQ8_63_19_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_19_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_158 = _weightQ8_63_19_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_19_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_159 = _weightQ8_63_19_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_19_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_160 = _weightQ8_63_19_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_19_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_161 = _weightQ8_63_19_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_19_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_162 = _weightQ8_63_19_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_19_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_163 = _weightQ8_63_19_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_19_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_164 = _weightQ8_63_19_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_19_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_165 = _weightQ8_63_19_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_19_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_166 = _weightQ8_63_19_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_19_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_167 = _weightQ8_63_19_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_19_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_168 = _weightQ8_63_19_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_19_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_169 = _weightQ8_63_19_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_19_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_170 = _weightQ8_63_19_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_19_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_171 = _weightQ8_63_19_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_19_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_172 = _weightQ8_63_19_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_19_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_173 = _weightQ8_63_19_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_19_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_174 = _weightQ8_63_19_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_19_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_175 = _weightQ8_63_19_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_19_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_176 = _weightQ8_63_19_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_19_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_177 = _weightQ8_63_19_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_19_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_178 = _weightQ8_63_19_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_19_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_179 = _weightQ8_63_19_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_19_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_180 = _weightQ8_63_19_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_19_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_181 = _weightQ8_63_19_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_19_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_182 = _weightQ8_63_19_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_19_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_183 = _weightQ8_63_19_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_19_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_184 = _weightQ8_63_19_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_19_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_185 = _weightQ8_63_19_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_19_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_186 = _weightQ8_63_19_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_19_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_187 = _weightQ8_63_19_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_19_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_188 = _weightQ8_63_19_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_19_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_leadingZeros_T_189 = _weightQ8_63_19_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_19_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_19_leadingZeros = _weightQ8_63_19_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_19_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_19_expRaw_T_1 = 6'h1f - weightQ8_63_19_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_19_expRaw = weightQ8_63_19_isZero ? 6'h0 : _weightQ8_63_19_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_19_shiftAmt_T_2 = weightQ8_63_19_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_19_shiftAmt = weightQ8_63_19_expRaw > 6'h3 ? _weightQ8_63_19_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_19_mantissaRaw_T = weightQ8_63_19_absClipped >> weightQ8_63_19_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_19_mantissaRaw = _weightQ8_63_19_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_19_mantissa = weightQ8_63_19_expRaw >= 6'h3 ? weightQ8_63_19_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_19_expAdjusted = weightQ8_63_19_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_19_exp_T_4 = weightQ8_63_19_expAdjusted > 7'hf ? 4'hf : weightQ8_63_19_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_19_exp = weightQ8_63_19_isZero ? 4'h0 : _weightQ8_63_19_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_19_fp8 = {weightQ8_63_19_clippedX[31],weightQ8_63_19_exp,weightQ8_63_19_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_20_T = {24'h0,linear_weight_63_20}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_20_sign = _weightQ8_63_20_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_20_absX_T = ~_weightQ8_63_20_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_20_absX_T_2 = _weightQ8_63_20_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_20_absX = weightQ8_63_20_sign ? _weightQ8_63_20_absX_T_2 : _weightQ8_63_20_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_20_shiftedX_T_1 = _GEN_14432 - weightQ8_63_20_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_20_shiftedX_T_3 = weightQ8_63_20_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_20_shiftedX = weightQ8_63_20_sign ? _weightQ8_63_20_shiftedX_T_1 :
    _weightQ8_63_20_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_20_scaledX_T_1 = weightQ8_63_20_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_20_scaledX = _weightQ8_63_20_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_20_clippedX_T_2 = weightQ8_63_20_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_20_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_20_clippedX = weightQ8_63_20_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_20_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_20_absClipped_T_1 = ~weightQ8_63_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_20_absClipped_T_3 = _weightQ8_63_20_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_20_absClipped = weightQ8_63_20_clippedX[31] ? _weightQ8_63_20_absClipped_T_3 :
    weightQ8_63_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_20_isZero = weightQ8_63_20_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37534 = {{16'd0}, weightQ8_63_20_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_4 = _GEN_37534 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_6 = {weightQ8_63_20_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_8 = _weightQ8_63_20_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_9 = _weightQ8_63_20_leadingZeros_T_4 | _weightQ8_63_20_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37535 = {{8'd0}, _weightQ8_63_20_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_14 = _GEN_37535 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_16 = {_weightQ8_63_20_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_18 = _weightQ8_63_20_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_19 = _weightQ8_63_20_leadingZeros_T_14 | _weightQ8_63_20_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37536 = {{4'd0}, _weightQ8_63_20_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_24 = _GEN_37536 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_26 = {_weightQ8_63_20_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_28 = _weightQ8_63_20_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_29 = _weightQ8_63_20_leadingZeros_T_24 | _weightQ8_63_20_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37537 = {{2'd0}, _weightQ8_63_20_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_34 = _GEN_37537 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_36 = {_weightQ8_63_20_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_38 = _weightQ8_63_20_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_39 = _weightQ8_63_20_leadingZeros_T_34 | _weightQ8_63_20_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37538 = {{1'd0}, _weightQ8_63_20_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_44 = _GEN_37538 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_46 = {_weightQ8_63_20_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_48 = _weightQ8_63_20_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_20_leadingZeros_T_49 = _weightQ8_63_20_leadingZeros_T_44 | _weightQ8_63_20_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37539 = {{8'd0}, weightQ8_63_20_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_55 = _GEN_37539 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_57 = {weightQ8_63_20_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_59 = _weightQ8_63_20_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_60 = _weightQ8_63_20_leadingZeros_T_55 | _weightQ8_63_20_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37540 = {{4'd0}, _weightQ8_63_20_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_65 = _GEN_37540 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_67 = {_weightQ8_63_20_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_69 = _weightQ8_63_20_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_70 = _weightQ8_63_20_leadingZeros_T_65 | _weightQ8_63_20_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37541 = {{2'd0}, _weightQ8_63_20_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_75 = _GEN_37541 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_77 = {_weightQ8_63_20_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_79 = _weightQ8_63_20_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_80 = _weightQ8_63_20_leadingZeros_T_75 | _weightQ8_63_20_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37542 = {{1'd0}, _weightQ8_63_20_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_85 = _GEN_37542 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_87 = {_weightQ8_63_20_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_89 = _weightQ8_63_20_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_20_leadingZeros_T_90 = _weightQ8_63_20_leadingZeros_T_85 | _weightQ8_63_20_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_20_leadingZeros_T_93 = {_weightQ8_63_20_leadingZeros_T_49,_weightQ8_63_20_leadingZeros_T_90,
    weightQ8_63_20_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_143 = _weightQ8_63_20_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_144 = _weightQ8_63_20_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_20_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_145 = _weightQ8_63_20_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_20_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_146 = _weightQ8_63_20_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_20_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_147 = _weightQ8_63_20_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_20_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_148 = _weightQ8_63_20_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_20_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_149 = _weightQ8_63_20_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_20_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_150 = _weightQ8_63_20_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_20_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_151 = _weightQ8_63_20_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_20_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_152 = _weightQ8_63_20_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_20_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_153 = _weightQ8_63_20_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_20_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_154 = _weightQ8_63_20_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_20_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_155 = _weightQ8_63_20_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_20_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_156 = _weightQ8_63_20_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_20_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_157 = _weightQ8_63_20_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_20_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_158 = _weightQ8_63_20_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_20_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_159 = _weightQ8_63_20_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_20_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_160 = _weightQ8_63_20_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_20_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_161 = _weightQ8_63_20_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_20_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_162 = _weightQ8_63_20_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_20_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_163 = _weightQ8_63_20_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_20_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_164 = _weightQ8_63_20_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_20_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_165 = _weightQ8_63_20_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_20_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_166 = _weightQ8_63_20_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_20_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_167 = _weightQ8_63_20_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_20_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_168 = _weightQ8_63_20_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_20_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_169 = _weightQ8_63_20_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_20_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_170 = _weightQ8_63_20_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_20_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_171 = _weightQ8_63_20_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_20_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_172 = _weightQ8_63_20_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_20_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_173 = _weightQ8_63_20_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_20_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_174 = _weightQ8_63_20_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_20_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_175 = _weightQ8_63_20_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_20_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_176 = _weightQ8_63_20_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_20_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_177 = _weightQ8_63_20_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_20_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_178 = _weightQ8_63_20_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_20_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_179 = _weightQ8_63_20_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_20_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_180 = _weightQ8_63_20_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_20_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_181 = _weightQ8_63_20_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_20_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_182 = _weightQ8_63_20_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_20_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_183 = _weightQ8_63_20_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_20_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_184 = _weightQ8_63_20_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_20_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_185 = _weightQ8_63_20_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_20_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_186 = _weightQ8_63_20_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_20_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_187 = _weightQ8_63_20_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_20_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_188 = _weightQ8_63_20_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_20_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_leadingZeros_T_189 = _weightQ8_63_20_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_20_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_20_leadingZeros = _weightQ8_63_20_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_20_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_20_expRaw_T_1 = 6'h1f - weightQ8_63_20_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_20_expRaw = weightQ8_63_20_isZero ? 6'h0 : _weightQ8_63_20_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_20_shiftAmt_T_2 = weightQ8_63_20_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_20_shiftAmt = weightQ8_63_20_expRaw > 6'h3 ? _weightQ8_63_20_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_20_mantissaRaw_T = weightQ8_63_20_absClipped >> weightQ8_63_20_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_20_mantissaRaw = _weightQ8_63_20_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_20_mantissa = weightQ8_63_20_expRaw >= 6'h3 ? weightQ8_63_20_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_20_expAdjusted = weightQ8_63_20_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_20_exp_T_4 = weightQ8_63_20_expAdjusted > 7'hf ? 4'hf : weightQ8_63_20_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_20_exp = weightQ8_63_20_isZero ? 4'h0 : _weightQ8_63_20_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_20_fp8 = {weightQ8_63_20_clippedX[31],weightQ8_63_20_exp,weightQ8_63_20_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_21_T = {24'h0,linear_weight_63_21}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_21_sign = _weightQ8_63_21_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_21_absX_T = ~_weightQ8_63_21_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_21_absX_T_2 = _weightQ8_63_21_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_21_absX = weightQ8_63_21_sign ? _weightQ8_63_21_absX_T_2 : _weightQ8_63_21_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_21_shiftedX_T_1 = _GEN_14432 - weightQ8_63_21_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_21_shiftedX_T_3 = weightQ8_63_21_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_21_shiftedX = weightQ8_63_21_sign ? _weightQ8_63_21_shiftedX_T_1 :
    _weightQ8_63_21_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_21_scaledX_T_1 = weightQ8_63_21_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_21_scaledX = _weightQ8_63_21_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_21_clippedX_T_2 = weightQ8_63_21_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_21_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_21_clippedX = weightQ8_63_21_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_21_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_21_absClipped_T_1 = ~weightQ8_63_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_21_absClipped_T_3 = _weightQ8_63_21_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_21_absClipped = weightQ8_63_21_clippedX[31] ? _weightQ8_63_21_absClipped_T_3 :
    weightQ8_63_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_21_isZero = weightQ8_63_21_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37545 = {{16'd0}, weightQ8_63_21_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_4 = _GEN_37545 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_6 = {weightQ8_63_21_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_8 = _weightQ8_63_21_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_9 = _weightQ8_63_21_leadingZeros_T_4 | _weightQ8_63_21_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37546 = {{8'd0}, _weightQ8_63_21_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_14 = _GEN_37546 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_16 = {_weightQ8_63_21_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_18 = _weightQ8_63_21_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_19 = _weightQ8_63_21_leadingZeros_T_14 | _weightQ8_63_21_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37547 = {{4'd0}, _weightQ8_63_21_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_24 = _GEN_37547 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_26 = {_weightQ8_63_21_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_28 = _weightQ8_63_21_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_29 = _weightQ8_63_21_leadingZeros_T_24 | _weightQ8_63_21_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37548 = {{2'd0}, _weightQ8_63_21_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_34 = _GEN_37548 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_36 = {_weightQ8_63_21_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_38 = _weightQ8_63_21_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_39 = _weightQ8_63_21_leadingZeros_T_34 | _weightQ8_63_21_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37549 = {{1'd0}, _weightQ8_63_21_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_44 = _GEN_37549 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_46 = {_weightQ8_63_21_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_48 = _weightQ8_63_21_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_21_leadingZeros_T_49 = _weightQ8_63_21_leadingZeros_T_44 | _weightQ8_63_21_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37550 = {{8'd0}, weightQ8_63_21_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_55 = _GEN_37550 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_57 = {weightQ8_63_21_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_59 = _weightQ8_63_21_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_60 = _weightQ8_63_21_leadingZeros_T_55 | _weightQ8_63_21_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37551 = {{4'd0}, _weightQ8_63_21_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_65 = _GEN_37551 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_67 = {_weightQ8_63_21_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_69 = _weightQ8_63_21_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_70 = _weightQ8_63_21_leadingZeros_T_65 | _weightQ8_63_21_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37552 = {{2'd0}, _weightQ8_63_21_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_75 = _GEN_37552 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_77 = {_weightQ8_63_21_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_79 = _weightQ8_63_21_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_80 = _weightQ8_63_21_leadingZeros_T_75 | _weightQ8_63_21_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37553 = {{1'd0}, _weightQ8_63_21_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_85 = _GEN_37553 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_87 = {_weightQ8_63_21_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_89 = _weightQ8_63_21_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_21_leadingZeros_T_90 = _weightQ8_63_21_leadingZeros_T_85 | _weightQ8_63_21_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_21_leadingZeros_T_93 = {_weightQ8_63_21_leadingZeros_T_49,_weightQ8_63_21_leadingZeros_T_90,
    weightQ8_63_21_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_143 = _weightQ8_63_21_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_144 = _weightQ8_63_21_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_21_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_145 = _weightQ8_63_21_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_21_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_146 = _weightQ8_63_21_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_21_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_147 = _weightQ8_63_21_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_21_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_148 = _weightQ8_63_21_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_21_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_149 = _weightQ8_63_21_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_21_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_150 = _weightQ8_63_21_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_21_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_151 = _weightQ8_63_21_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_21_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_152 = _weightQ8_63_21_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_21_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_153 = _weightQ8_63_21_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_21_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_154 = _weightQ8_63_21_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_21_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_155 = _weightQ8_63_21_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_21_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_156 = _weightQ8_63_21_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_21_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_157 = _weightQ8_63_21_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_21_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_158 = _weightQ8_63_21_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_21_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_159 = _weightQ8_63_21_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_21_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_160 = _weightQ8_63_21_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_21_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_161 = _weightQ8_63_21_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_21_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_162 = _weightQ8_63_21_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_21_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_163 = _weightQ8_63_21_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_21_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_164 = _weightQ8_63_21_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_21_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_165 = _weightQ8_63_21_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_21_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_166 = _weightQ8_63_21_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_21_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_167 = _weightQ8_63_21_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_21_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_168 = _weightQ8_63_21_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_21_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_169 = _weightQ8_63_21_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_21_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_170 = _weightQ8_63_21_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_21_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_171 = _weightQ8_63_21_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_21_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_172 = _weightQ8_63_21_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_21_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_173 = _weightQ8_63_21_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_21_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_174 = _weightQ8_63_21_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_21_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_175 = _weightQ8_63_21_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_21_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_176 = _weightQ8_63_21_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_21_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_177 = _weightQ8_63_21_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_21_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_178 = _weightQ8_63_21_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_21_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_179 = _weightQ8_63_21_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_21_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_180 = _weightQ8_63_21_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_21_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_181 = _weightQ8_63_21_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_21_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_182 = _weightQ8_63_21_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_21_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_183 = _weightQ8_63_21_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_21_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_184 = _weightQ8_63_21_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_21_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_185 = _weightQ8_63_21_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_21_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_186 = _weightQ8_63_21_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_21_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_187 = _weightQ8_63_21_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_21_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_188 = _weightQ8_63_21_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_21_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_leadingZeros_T_189 = _weightQ8_63_21_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_21_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_21_leadingZeros = _weightQ8_63_21_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_21_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_21_expRaw_T_1 = 6'h1f - weightQ8_63_21_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_21_expRaw = weightQ8_63_21_isZero ? 6'h0 : _weightQ8_63_21_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_21_shiftAmt_T_2 = weightQ8_63_21_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_21_shiftAmt = weightQ8_63_21_expRaw > 6'h3 ? _weightQ8_63_21_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_21_mantissaRaw_T = weightQ8_63_21_absClipped >> weightQ8_63_21_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_21_mantissaRaw = _weightQ8_63_21_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_21_mantissa = weightQ8_63_21_expRaw >= 6'h3 ? weightQ8_63_21_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_21_expAdjusted = weightQ8_63_21_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_21_exp_T_4 = weightQ8_63_21_expAdjusted > 7'hf ? 4'hf : weightQ8_63_21_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_21_exp = weightQ8_63_21_isZero ? 4'h0 : _weightQ8_63_21_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_21_fp8 = {weightQ8_63_21_clippedX[31],weightQ8_63_21_exp,weightQ8_63_21_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_22_T = {24'h0,linear_weight_63_22}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_22_sign = _weightQ8_63_22_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_22_absX_T = ~_weightQ8_63_22_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_22_absX_T_2 = _weightQ8_63_22_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_22_absX = weightQ8_63_22_sign ? _weightQ8_63_22_absX_T_2 : _weightQ8_63_22_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_22_shiftedX_T_1 = _GEN_14432 - weightQ8_63_22_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_22_shiftedX_T_3 = weightQ8_63_22_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_22_shiftedX = weightQ8_63_22_sign ? _weightQ8_63_22_shiftedX_T_1 :
    _weightQ8_63_22_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_22_scaledX_T_1 = weightQ8_63_22_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_22_scaledX = _weightQ8_63_22_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_22_clippedX_T_2 = weightQ8_63_22_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_22_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_22_clippedX = weightQ8_63_22_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_22_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_22_absClipped_T_1 = ~weightQ8_63_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_22_absClipped_T_3 = _weightQ8_63_22_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_22_absClipped = weightQ8_63_22_clippedX[31] ? _weightQ8_63_22_absClipped_T_3 :
    weightQ8_63_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_22_isZero = weightQ8_63_22_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37556 = {{16'd0}, weightQ8_63_22_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_4 = _GEN_37556 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_6 = {weightQ8_63_22_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_8 = _weightQ8_63_22_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_9 = _weightQ8_63_22_leadingZeros_T_4 | _weightQ8_63_22_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37557 = {{8'd0}, _weightQ8_63_22_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_14 = _GEN_37557 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_16 = {_weightQ8_63_22_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_18 = _weightQ8_63_22_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_19 = _weightQ8_63_22_leadingZeros_T_14 | _weightQ8_63_22_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37558 = {{4'd0}, _weightQ8_63_22_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_24 = _GEN_37558 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_26 = {_weightQ8_63_22_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_28 = _weightQ8_63_22_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_29 = _weightQ8_63_22_leadingZeros_T_24 | _weightQ8_63_22_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37559 = {{2'd0}, _weightQ8_63_22_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_34 = _GEN_37559 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_36 = {_weightQ8_63_22_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_38 = _weightQ8_63_22_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_39 = _weightQ8_63_22_leadingZeros_T_34 | _weightQ8_63_22_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37560 = {{1'd0}, _weightQ8_63_22_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_44 = _GEN_37560 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_46 = {_weightQ8_63_22_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_48 = _weightQ8_63_22_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_22_leadingZeros_T_49 = _weightQ8_63_22_leadingZeros_T_44 | _weightQ8_63_22_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37561 = {{8'd0}, weightQ8_63_22_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_55 = _GEN_37561 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_57 = {weightQ8_63_22_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_59 = _weightQ8_63_22_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_60 = _weightQ8_63_22_leadingZeros_T_55 | _weightQ8_63_22_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37562 = {{4'd0}, _weightQ8_63_22_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_65 = _GEN_37562 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_67 = {_weightQ8_63_22_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_69 = _weightQ8_63_22_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_70 = _weightQ8_63_22_leadingZeros_T_65 | _weightQ8_63_22_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37563 = {{2'd0}, _weightQ8_63_22_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_75 = _GEN_37563 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_77 = {_weightQ8_63_22_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_79 = _weightQ8_63_22_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_80 = _weightQ8_63_22_leadingZeros_T_75 | _weightQ8_63_22_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37564 = {{1'd0}, _weightQ8_63_22_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_85 = _GEN_37564 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_87 = {_weightQ8_63_22_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_89 = _weightQ8_63_22_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_22_leadingZeros_T_90 = _weightQ8_63_22_leadingZeros_T_85 | _weightQ8_63_22_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_22_leadingZeros_T_93 = {_weightQ8_63_22_leadingZeros_T_49,_weightQ8_63_22_leadingZeros_T_90,
    weightQ8_63_22_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_143 = _weightQ8_63_22_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_144 = _weightQ8_63_22_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_22_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_145 = _weightQ8_63_22_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_22_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_146 = _weightQ8_63_22_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_22_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_147 = _weightQ8_63_22_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_22_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_148 = _weightQ8_63_22_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_22_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_149 = _weightQ8_63_22_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_22_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_150 = _weightQ8_63_22_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_22_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_151 = _weightQ8_63_22_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_22_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_152 = _weightQ8_63_22_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_22_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_153 = _weightQ8_63_22_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_22_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_154 = _weightQ8_63_22_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_22_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_155 = _weightQ8_63_22_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_22_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_156 = _weightQ8_63_22_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_22_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_157 = _weightQ8_63_22_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_22_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_158 = _weightQ8_63_22_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_22_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_159 = _weightQ8_63_22_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_22_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_160 = _weightQ8_63_22_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_22_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_161 = _weightQ8_63_22_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_22_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_162 = _weightQ8_63_22_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_22_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_163 = _weightQ8_63_22_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_22_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_164 = _weightQ8_63_22_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_22_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_165 = _weightQ8_63_22_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_22_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_166 = _weightQ8_63_22_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_22_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_167 = _weightQ8_63_22_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_22_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_168 = _weightQ8_63_22_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_22_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_169 = _weightQ8_63_22_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_22_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_170 = _weightQ8_63_22_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_22_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_171 = _weightQ8_63_22_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_22_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_172 = _weightQ8_63_22_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_22_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_173 = _weightQ8_63_22_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_22_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_174 = _weightQ8_63_22_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_22_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_175 = _weightQ8_63_22_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_22_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_176 = _weightQ8_63_22_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_22_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_177 = _weightQ8_63_22_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_22_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_178 = _weightQ8_63_22_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_22_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_179 = _weightQ8_63_22_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_22_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_180 = _weightQ8_63_22_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_22_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_181 = _weightQ8_63_22_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_22_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_182 = _weightQ8_63_22_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_22_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_183 = _weightQ8_63_22_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_22_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_184 = _weightQ8_63_22_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_22_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_185 = _weightQ8_63_22_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_22_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_186 = _weightQ8_63_22_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_22_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_187 = _weightQ8_63_22_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_22_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_188 = _weightQ8_63_22_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_22_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_leadingZeros_T_189 = _weightQ8_63_22_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_22_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_22_leadingZeros = _weightQ8_63_22_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_22_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_22_expRaw_T_1 = 6'h1f - weightQ8_63_22_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_22_expRaw = weightQ8_63_22_isZero ? 6'h0 : _weightQ8_63_22_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_22_shiftAmt_T_2 = weightQ8_63_22_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_22_shiftAmt = weightQ8_63_22_expRaw > 6'h3 ? _weightQ8_63_22_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_22_mantissaRaw_T = weightQ8_63_22_absClipped >> weightQ8_63_22_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_22_mantissaRaw = _weightQ8_63_22_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_22_mantissa = weightQ8_63_22_expRaw >= 6'h3 ? weightQ8_63_22_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_22_expAdjusted = weightQ8_63_22_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_22_exp_T_4 = weightQ8_63_22_expAdjusted > 7'hf ? 4'hf : weightQ8_63_22_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_22_exp = weightQ8_63_22_isZero ? 4'h0 : _weightQ8_63_22_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_22_fp8 = {weightQ8_63_22_clippedX[31],weightQ8_63_22_exp,weightQ8_63_22_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_23_T = {24'h0,linear_weight_63_23}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_23_sign = _weightQ8_63_23_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_23_absX_T = ~_weightQ8_63_23_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_23_absX_T_2 = _weightQ8_63_23_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_23_absX = weightQ8_63_23_sign ? _weightQ8_63_23_absX_T_2 : _weightQ8_63_23_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_23_shiftedX_T_1 = _GEN_14432 - weightQ8_63_23_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_23_shiftedX_T_3 = weightQ8_63_23_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_23_shiftedX = weightQ8_63_23_sign ? _weightQ8_63_23_shiftedX_T_1 :
    _weightQ8_63_23_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_23_scaledX_T_1 = weightQ8_63_23_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_23_scaledX = _weightQ8_63_23_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_23_clippedX_T_2 = weightQ8_63_23_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_23_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_23_clippedX = weightQ8_63_23_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_23_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_23_absClipped_T_1 = ~weightQ8_63_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_23_absClipped_T_3 = _weightQ8_63_23_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_23_absClipped = weightQ8_63_23_clippedX[31] ? _weightQ8_63_23_absClipped_T_3 :
    weightQ8_63_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_23_isZero = weightQ8_63_23_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37567 = {{16'd0}, weightQ8_63_23_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_4 = _GEN_37567 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_6 = {weightQ8_63_23_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_8 = _weightQ8_63_23_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_9 = _weightQ8_63_23_leadingZeros_T_4 | _weightQ8_63_23_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37568 = {{8'd0}, _weightQ8_63_23_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_14 = _GEN_37568 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_16 = {_weightQ8_63_23_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_18 = _weightQ8_63_23_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_19 = _weightQ8_63_23_leadingZeros_T_14 | _weightQ8_63_23_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37569 = {{4'd0}, _weightQ8_63_23_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_24 = _GEN_37569 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_26 = {_weightQ8_63_23_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_28 = _weightQ8_63_23_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_29 = _weightQ8_63_23_leadingZeros_T_24 | _weightQ8_63_23_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37570 = {{2'd0}, _weightQ8_63_23_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_34 = _GEN_37570 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_36 = {_weightQ8_63_23_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_38 = _weightQ8_63_23_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_39 = _weightQ8_63_23_leadingZeros_T_34 | _weightQ8_63_23_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37571 = {{1'd0}, _weightQ8_63_23_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_44 = _GEN_37571 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_46 = {_weightQ8_63_23_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_48 = _weightQ8_63_23_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_23_leadingZeros_T_49 = _weightQ8_63_23_leadingZeros_T_44 | _weightQ8_63_23_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37572 = {{8'd0}, weightQ8_63_23_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_55 = _GEN_37572 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_57 = {weightQ8_63_23_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_59 = _weightQ8_63_23_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_60 = _weightQ8_63_23_leadingZeros_T_55 | _weightQ8_63_23_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37573 = {{4'd0}, _weightQ8_63_23_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_65 = _GEN_37573 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_67 = {_weightQ8_63_23_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_69 = _weightQ8_63_23_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_70 = _weightQ8_63_23_leadingZeros_T_65 | _weightQ8_63_23_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37574 = {{2'd0}, _weightQ8_63_23_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_75 = _GEN_37574 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_77 = {_weightQ8_63_23_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_79 = _weightQ8_63_23_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_80 = _weightQ8_63_23_leadingZeros_T_75 | _weightQ8_63_23_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37575 = {{1'd0}, _weightQ8_63_23_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_85 = _GEN_37575 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_87 = {_weightQ8_63_23_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_89 = _weightQ8_63_23_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_23_leadingZeros_T_90 = _weightQ8_63_23_leadingZeros_T_85 | _weightQ8_63_23_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_23_leadingZeros_T_93 = {_weightQ8_63_23_leadingZeros_T_49,_weightQ8_63_23_leadingZeros_T_90,
    weightQ8_63_23_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_143 = _weightQ8_63_23_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_144 = _weightQ8_63_23_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_23_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_145 = _weightQ8_63_23_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_23_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_146 = _weightQ8_63_23_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_23_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_147 = _weightQ8_63_23_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_23_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_148 = _weightQ8_63_23_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_23_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_149 = _weightQ8_63_23_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_23_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_150 = _weightQ8_63_23_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_23_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_151 = _weightQ8_63_23_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_23_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_152 = _weightQ8_63_23_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_23_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_153 = _weightQ8_63_23_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_23_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_154 = _weightQ8_63_23_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_23_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_155 = _weightQ8_63_23_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_23_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_156 = _weightQ8_63_23_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_23_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_157 = _weightQ8_63_23_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_23_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_158 = _weightQ8_63_23_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_23_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_159 = _weightQ8_63_23_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_23_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_160 = _weightQ8_63_23_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_23_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_161 = _weightQ8_63_23_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_23_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_162 = _weightQ8_63_23_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_23_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_163 = _weightQ8_63_23_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_23_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_164 = _weightQ8_63_23_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_23_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_165 = _weightQ8_63_23_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_23_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_166 = _weightQ8_63_23_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_23_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_167 = _weightQ8_63_23_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_23_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_168 = _weightQ8_63_23_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_23_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_169 = _weightQ8_63_23_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_23_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_170 = _weightQ8_63_23_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_23_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_171 = _weightQ8_63_23_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_23_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_172 = _weightQ8_63_23_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_23_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_173 = _weightQ8_63_23_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_23_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_174 = _weightQ8_63_23_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_23_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_175 = _weightQ8_63_23_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_23_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_176 = _weightQ8_63_23_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_23_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_177 = _weightQ8_63_23_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_23_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_178 = _weightQ8_63_23_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_23_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_179 = _weightQ8_63_23_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_23_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_180 = _weightQ8_63_23_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_23_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_181 = _weightQ8_63_23_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_23_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_182 = _weightQ8_63_23_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_23_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_183 = _weightQ8_63_23_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_23_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_184 = _weightQ8_63_23_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_23_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_185 = _weightQ8_63_23_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_23_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_186 = _weightQ8_63_23_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_23_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_187 = _weightQ8_63_23_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_23_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_188 = _weightQ8_63_23_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_23_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_leadingZeros_T_189 = _weightQ8_63_23_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_23_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_23_leadingZeros = _weightQ8_63_23_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_23_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_23_expRaw_T_1 = 6'h1f - weightQ8_63_23_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_23_expRaw = weightQ8_63_23_isZero ? 6'h0 : _weightQ8_63_23_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_23_shiftAmt_T_2 = weightQ8_63_23_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_23_shiftAmt = weightQ8_63_23_expRaw > 6'h3 ? _weightQ8_63_23_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_23_mantissaRaw_T = weightQ8_63_23_absClipped >> weightQ8_63_23_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_23_mantissaRaw = _weightQ8_63_23_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_23_mantissa = weightQ8_63_23_expRaw >= 6'h3 ? weightQ8_63_23_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_23_expAdjusted = weightQ8_63_23_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_23_exp_T_4 = weightQ8_63_23_expAdjusted > 7'hf ? 4'hf : weightQ8_63_23_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_23_exp = weightQ8_63_23_isZero ? 4'h0 : _weightQ8_63_23_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_23_fp8 = {weightQ8_63_23_clippedX[31],weightQ8_63_23_exp,weightQ8_63_23_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_24_T = {24'h0,linear_weight_63_24}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_24_sign = _weightQ8_63_24_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_24_absX_T = ~_weightQ8_63_24_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_24_absX_T_2 = _weightQ8_63_24_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_24_absX = weightQ8_63_24_sign ? _weightQ8_63_24_absX_T_2 : _weightQ8_63_24_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_24_shiftedX_T_1 = _GEN_14432 - weightQ8_63_24_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_24_shiftedX_T_3 = weightQ8_63_24_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_24_shiftedX = weightQ8_63_24_sign ? _weightQ8_63_24_shiftedX_T_1 :
    _weightQ8_63_24_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_24_scaledX_T_1 = weightQ8_63_24_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_24_scaledX = _weightQ8_63_24_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_24_clippedX_T_2 = weightQ8_63_24_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_24_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_24_clippedX = weightQ8_63_24_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_24_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_24_absClipped_T_1 = ~weightQ8_63_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_24_absClipped_T_3 = _weightQ8_63_24_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_24_absClipped = weightQ8_63_24_clippedX[31] ? _weightQ8_63_24_absClipped_T_3 :
    weightQ8_63_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_24_isZero = weightQ8_63_24_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37578 = {{16'd0}, weightQ8_63_24_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_4 = _GEN_37578 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_6 = {weightQ8_63_24_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_8 = _weightQ8_63_24_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_9 = _weightQ8_63_24_leadingZeros_T_4 | _weightQ8_63_24_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37579 = {{8'd0}, _weightQ8_63_24_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_14 = _GEN_37579 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_16 = {_weightQ8_63_24_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_18 = _weightQ8_63_24_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_19 = _weightQ8_63_24_leadingZeros_T_14 | _weightQ8_63_24_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37580 = {{4'd0}, _weightQ8_63_24_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_24 = _GEN_37580 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_26 = {_weightQ8_63_24_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_28 = _weightQ8_63_24_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_29 = _weightQ8_63_24_leadingZeros_T_24 | _weightQ8_63_24_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37581 = {{2'd0}, _weightQ8_63_24_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_34 = _GEN_37581 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_36 = {_weightQ8_63_24_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_38 = _weightQ8_63_24_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_39 = _weightQ8_63_24_leadingZeros_T_34 | _weightQ8_63_24_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37582 = {{1'd0}, _weightQ8_63_24_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_44 = _GEN_37582 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_46 = {_weightQ8_63_24_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_48 = _weightQ8_63_24_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_24_leadingZeros_T_49 = _weightQ8_63_24_leadingZeros_T_44 | _weightQ8_63_24_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37583 = {{8'd0}, weightQ8_63_24_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_55 = _GEN_37583 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_57 = {weightQ8_63_24_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_59 = _weightQ8_63_24_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_60 = _weightQ8_63_24_leadingZeros_T_55 | _weightQ8_63_24_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37584 = {{4'd0}, _weightQ8_63_24_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_65 = _GEN_37584 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_67 = {_weightQ8_63_24_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_69 = _weightQ8_63_24_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_70 = _weightQ8_63_24_leadingZeros_T_65 | _weightQ8_63_24_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37585 = {{2'd0}, _weightQ8_63_24_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_75 = _GEN_37585 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_77 = {_weightQ8_63_24_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_79 = _weightQ8_63_24_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_80 = _weightQ8_63_24_leadingZeros_T_75 | _weightQ8_63_24_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37586 = {{1'd0}, _weightQ8_63_24_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_85 = _GEN_37586 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_87 = {_weightQ8_63_24_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_89 = _weightQ8_63_24_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_24_leadingZeros_T_90 = _weightQ8_63_24_leadingZeros_T_85 | _weightQ8_63_24_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_24_leadingZeros_T_93 = {_weightQ8_63_24_leadingZeros_T_49,_weightQ8_63_24_leadingZeros_T_90,
    weightQ8_63_24_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_143 = _weightQ8_63_24_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_144 = _weightQ8_63_24_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_24_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_145 = _weightQ8_63_24_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_24_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_146 = _weightQ8_63_24_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_24_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_147 = _weightQ8_63_24_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_24_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_148 = _weightQ8_63_24_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_24_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_149 = _weightQ8_63_24_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_24_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_150 = _weightQ8_63_24_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_24_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_151 = _weightQ8_63_24_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_24_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_152 = _weightQ8_63_24_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_24_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_153 = _weightQ8_63_24_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_24_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_154 = _weightQ8_63_24_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_24_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_155 = _weightQ8_63_24_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_24_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_156 = _weightQ8_63_24_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_24_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_157 = _weightQ8_63_24_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_24_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_158 = _weightQ8_63_24_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_24_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_159 = _weightQ8_63_24_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_24_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_160 = _weightQ8_63_24_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_24_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_161 = _weightQ8_63_24_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_24_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_162 = _weightQ8_63_24_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_24_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_163 = _weightQ8_63_24_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_24_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_164 = _weightQ8_63_24_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_24_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_165 = _weightQ8_63_24_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_24_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_166 = _weightQ8_63_24_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_24_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_167 = _weightQ8_63_24_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_24_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_168 = _weightQ8_63_24_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_24_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_169 = _weightQ8_63_24_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_24_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_170 = _weightQ8_63_24_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_24_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_171 = _weightQ8_63_24_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_24_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_172 = _weightQ8_63_24_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_24_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_173 = _weightQ8_63_24_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_24_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_174 = _weightQ8_63_24_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_24_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_175 = _weightQ8_63_24_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_24_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_176 = _weightQ8_63_24_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_24_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_177 = _weightQ8_63_24_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_24_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_178 = _weightQ8_63_24_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_24_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_179 = _weightQ8_63_24_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_24_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_180 = _weightQ8_63_24_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_24_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_181 = _weightQ8_63_24_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_24_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_182 = _weightQ8_63_24_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_24_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_183 = _weightQ8_63_24_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_24_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_184 = _weightQ8_63_24_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_24_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_185 = _weightQ8_63_24_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_24_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_186 = _weightQ8_63_24_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_24_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_187 = _weightQ8_63_24_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_24_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_188 = _weightQ8_63_24_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_24_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_leadingZeros_T_189 = _weightQ8_63_24_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_24_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_24_leadingZeros = _weightQ8_63_24_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_24_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_24_expRaw_T_1 = 6'h1f - weightQ8_63_24_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_24_expRaw = weightQ8_63_24_isZero ? 6'h0 : _weightQ8_63_24_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_24_shiftAmt_T_2 = weightQ8_63_24_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_24_shiftAmt = weightQ8_63_24_expRaw > 6'h3 ? _weightQ8_63_24_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_24_mantissaRaw_T = weightQ8_63_24_absClipped >> weightQ8_63_24_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_24_mantissaRaw = _weightQ8_63_24_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_24_mantissa = weightQ8_63_24_expRaw >= 6'h3 ? weightQ8_63_24_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_24_expAdjusted = weightQ8_63_24_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_24_exp_T_4 = weightQ8_63_24_expAdjusted > 7'hf ? 4'hf : weightQ8_63_24_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_24_exp = weightQ8_63_24_isZero ? 4'h0 : _weightQ8_63_24_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_24_fp8 = {weightQ8_63_24_clippedX[31],weightQ8_63_24_exp,weightQ8_63_24_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_25_T = {24'h0,linear_weight_63_25}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_25_sign = _weightQ8_63_25_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_25_absX_T = ~_weightQ8_63_25_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_25_absX_T_2 = _weightQ8_63_25_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_25_absX = weightQ8_63_25_sign ? _weightQ8_63_25_absX_T_2 : _weightQ8_63_25_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_25_shiftedX_T_1 = _GEN_14432 - weightQ8_63_25_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_25_shiftedX_T_3 = weightQ8_63_25_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_25_shiftedX = weightQ8_63_25_sign ? _weightQ8_63_25_shiftedX_T_1 :
    _weightQ8_63_25_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_25_scaledX_T_1 = weightQ8_63_25_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_25_scaledX = _weightQ8_63_25_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_25_clippedX_T_2 = weightQ8_63_25_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_25_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_25_clippedX = weightQ8_63_25_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_25_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_25_absClipped_T_1 = ~weightQ8_63_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_25_absClipped_T_3 = _weightQ8_63_25_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_25_absClipped = weightQ8_63_25_clippedX[31] ? _weightQ8_63_25_absClipped_T_3 :
    weightQ8_63_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_25_isZero = weightQ8_63_25_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37589 = {{16'd0}, weightQ8_63_25_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_4 = _GEN_37589 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_6 = {weightQ8_63_25_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_8 = _weightQ8_63_25_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_9 = _weightQ8_63_25_leadingZeros_T_4 | _weightQ8_63_25_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37590 = {{8'd0}, _weightQ8_63_25_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_14 = _GEN_37590 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_16 = {_weightQ8_63_25_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_18 = _weightQ8_63_25_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_19 = _weightQ8_63_25_leadingZeros_T_14 | _weightQ8_63_25_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37591 = {{4'd0}, _weightQ8_63_25_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_24 = _GEN_37591 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_26 = {_weightQ8_63_25_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_28 = _weightQ8_63_25_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_29 = _weightQ8_63_25_leadingZeros_T_24 | _weightQ8_63_25_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37592 = {{2'd0}, _weightQ8_63_25_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_34 = _GEN_37592 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_36 = {_weightQ8_63_25_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_38 = _weightQ8_63_25_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_39 = _weightQ8_63_25_leadingZeros_T_34 | _weightQ8_63_25_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37593 = {{1'd0}, _weightQ8_63_25_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_44 = _GEN_37593 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_46 = {_weightQ8_63_25_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_48 = _weightQ8_63_25_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_25_leadingZeros_T_49 = _weightQ8_63_25_leadingZeros_T_44 | _weightQ8_63_25_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37594 = {{8'd0}, weightQ8_63_25_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_55 = _GEN_37594 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_57 = {weightQ8_63_25_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_59 = _weightQ8_63_25_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_60 = _weightQ8_63_25_leadingZeros_T_55 | _weightQ8_63_25_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37595 = {{4'd0}, _weightQ8_63_25_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_65 = _GEN_37595 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_67 = {_weightQ8_63_25_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_69 = _weightQ8_63_25_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_70 = _weightQ8_63_25_leadingZeros_T_65 | _weightQ8_63_25_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37596 = {{2'd0}, _weightQ8_63_25_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_75 = _GEN_37596 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_77 = {_weightQ8_63_25_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_79 = _weightQ8_63_25_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_80 = _weightQ8_63_25_leadingZeros_T_75 | _weightQ8_63_25_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37597 = {{1'd0}, _weightQ8_63_25_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_85 = _GEN_37597 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_87 = {_weightQ8_63_25_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_89 = _weightQ8_63_25_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_25_leadingZeros_T_90 = _weightQ8_63_25_leadingZeros_T_85 | _weightQ8_63_25_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_25_leadingZeros_T_93 = {_weightQ8_63_25_leadingZeros_T_49,_weightQ8_63_25_leadingZeros_T_90,
    weightQ8_63_25_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_143 = _weightQ8_63_25_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_144 = _weightQ8_63_25_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_25_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_145 = _weightQ8_63_25_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_25_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_146 = _weightQ8_63_25_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_25_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_147 = _weightQ8_63_25_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_25_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_148 = _weightQ8_63_25_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_25_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_149 = _weightQ8_63_25_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_25_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_150 = _weightQ8_63_25_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_25_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_151 = _weightQ8_63_25_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_25_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_152 = _weightQ8_63_25_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_25_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_153 = _weightQ8_63_25_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_25_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_154 = _weightQ8_63_25_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_25_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_155 = _weightQ8_63_25_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_25_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_156 = _weightQ8_63_25_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_25_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_157 = _weightQ8_63_25_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_25_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_158 = _weightQ8_63_25_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_25_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_159 = _weightQ8_63_25_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_25_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_160 = _weightQ8_63_25_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_25_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_161 = _weightQ8_63_25_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_25_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_162 = _weightQ8_63_25_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_25_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_163 = _weightQ8_63_25_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_25_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_164 = _weightQ8_63_25_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_25_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_165 = _weightQ8_63_25_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_25_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_166 = _weightQ8_63_25_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_25_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_167 = _weightQ8_63_25_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_25_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_168 = _weightQ8_63_25_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_25_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_169 = _weightQ8_63_25_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_25_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_170 = _weightQ8_63_25_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_25_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_171 = _weightQ8_63_25_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_25_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_172 = _weightQ8_63_25_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_25_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_173 = _weightQ8_63_25_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_25_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_174 = _weightQ8_63_25_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_25_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_175 = _weightQ8_63_25_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_25_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_176 = _weightQ8_63_25_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_25_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_177 = _weightQ8_63_25_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_25_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_178 = _weightQ8_63_25_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_25_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_179 = _weightQ8_63_25_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_25_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_180 = _weightQ8_63_25_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_25_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_181 = _weightQ8_63_25_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_25_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_182 = _weightQ8_63_25_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_25_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_183 = _weightQ8_63_25_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_25_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_184 = _weightQ8_63_25_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_25_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_185 = _weightQ8_63_25_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_25_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_186 = _weightQ8_63_25_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_25_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_187 = _weightQ8_63_25_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_25_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_188 = _weightQ8_63_25_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_25_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_leadingZeros_T_189 = _weightQ8_63_25_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_25_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_25_leadingZeros = _weightQ8_63_25_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_25_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_25_expRaw_T_1 = 6'h1f - weightQ8_63_25_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_25_expRaw = weightQ8_63_25_isZero ? 6'h0 : _weightQ8_63_25_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_25_shiftAmt_T_2 = weightQ8_63_25_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_25_shiftAmt = weightQ8_63_25_expRaw > 6'h3 ? _weightQ8_63_25_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_25_mantissaRaw_T = weightQ8_63_25_absClipped >> weightQ8_63_25_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_25_mantissaRaw = _weightQ8_63_25_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_25_mantissa = weightQ8_63_25_expRaw >= 6'h3 ? weightQ8_63_25_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_25_expAdjusted = weightQ8_63_25_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_25_exp_T_4 = weightQ8_63_25_expAdjusted > 7'hf ? 4'hf : weightQ8_63_25_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_25_exp = weightQ8_63_25_isZero ? 4'h0 : _weightQ8_63_25_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_25_fp8 = {weightQ8_63_25_clippedX[31],weightQ8_63_25_exp,weightQ8_63_25_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_26_T = {24'h0,linear_weight_63_26}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_26_sign = _weightQ8_63_26_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_26_absX_T = ~_weightQ8_63_26_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_26_absX_T_2 = _weightQ8_63_26_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_26_absX = weightQ8_63_26_sign ? _weightQ8_63_26_absX_T_2 : _weightQ8_63_26_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_26_shiftedX_T_1 = _GEN_14432 - weightQ8_63_26_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_26_shiftedX_T_3 = weightQ8_63_26_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_26_shiftedX = weightQ8_63_26_sign ? _weightQ8_63_26_shiftedX_T_1 :
    _weightQ8_63_26_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_26_scaledX_T_1 = weightQ8_63_26_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_26_scaledX = _weightQ8_63_26_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_26_clippedX_T_2 = weightQ8_63_26_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_26_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_26_clippedX = weightQ8_63_26_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_26_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_26_absClipped_T_1 = ~weightQ8_63_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_26_absClipped_T_3 = _weightQ8_63_26_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_26_absClipped = weightQ8_63_26_clippedX[31] ? _weightQ8_63_26_absClipped_T_3 :
    weightQ8_63_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_26_isZero = weightQ8_63_26_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37600 = {{16'd0}, weightQ8_63_26_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_4 = _GEN_37600 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_6 = {weightQ8_63_26_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_8 = _weightQ8_63_26_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_9 = _weightQ8_63_26_leadingZeros_T_4 | _weightQ8_63_26_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37601 = {{8'd0}, _weightQ8_63_26_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_14 = _GEN_37601 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_16 = {_weightQ8_63_26_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_18 = _weightQ8_63_26_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_19 = _weightQ8_63_26_leadingZeros_T_14 | _weightQ8_63_26_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37602 = {{4'd0}, _weightQ8_63_26_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_24 = _GEN_37602 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_26 = {_weightQ8_63_26_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_28 = _weightQ8_63_26_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_29 = _weightQ8_63_26_leadingZeros_T_24 | _weightQ8_63_26_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37603 = {{2'd0}, _weightQ8_63_26_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_34 = _GEN_37603 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_36 = {_weightQ8_63_26_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_38 = _weightQ8_63_26_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_39 = _weightQ8_63_26_leadingZeros_T_34 | _weightQ8_63_26_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37604 = {{1'd0}, _weightQ8_63_26_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_44 = _GEN_37604 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_46 = {_weightQ8_63_26_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_48 = _weightQ8_63_26_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_26_leadingZeros_T_49 = _weightQ8_63_26_leadingZeros_T_44 | _weightQ8_63_26_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37605 = {{8'd0}, weightQ8_63_26_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_55 = _GEN_37605 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_57 = {weightQ8_63_26_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_59 = _weightQ8_63_26_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_60 = _weightQ8_63_26_leadingZeros_T_55 | _weightQ8_63_26_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37606 = {{4'd0}, _weightQ8_63_26_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_65 = _GEN_37606 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_67 = {_weightQ8_63_26_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_69 = _weightQ8_63_26_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_70 = _weightQ8_63_26_leadingZeros_T_65 | _weightQ8_63_26_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37607 = {{2'd0}, _weightQ8_63_26_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_75 = _GEN_37607 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_77 = {_weightQ8_63_26_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_79 = _weightQ8_63_26_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_80 = _weightQ8_63_26_leadingZeros_T_75 | _weightQ8_63_26_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37608 = {{1'd0}, _weightQ8_63_26_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_85 = _GEN_37608 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_87 = {_weightQ8_63_26_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_89 = _weightQ8_63_26_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_26_leadingZeros_T_90 = _weightQ8_63_26_leadingZeros_T_85 | _weightQ8_63_26_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_26_leadingZeros_T_93 = {_weightQ8_63_26_leadingZeros_T_49,_weightQ8_63_26_leadingZeros_T_90,
    weightQ8_63_26_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_143 = _weightQ8_63_26_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_144 = _weightQ8_63_26_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_26_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_145 = _weightQ8_63_26_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_26_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_146 = _weightQ8_63_26_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_26_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_147 = _weightQ8_63_26_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_26_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_148 = _weightQ8_63_26_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_26_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_149 = _weightQ8_63_26_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_26_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_150 = _weightQ8_63_26_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_26_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_151 = _weightQ8_63_26_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_26_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_152 = _weightQ8_63_26_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_26_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_153 = _weightQ8_63_26_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_26_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_154 = _weightQ8_63_26_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_26_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_155 = _weightQ8_63_26_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_26_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_156 = _weightQ8_63_26_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_26_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_157 = _weightQ8_63_26_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_26_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_158 = _weightQ8_63_26_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_26_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_159 = _weightQ8_63_26_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_26_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_160 = _weightQ8_63_26_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_26_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_161 = _weightQ8_63_26_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_26_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_162 = _weightQ8_63_26_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_26_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_163 = _weightQ8_63_26_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_26_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_164 = _weightQ8_63_26_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_26_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_165 = _weightQ8_63_26_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_26_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_166 = _weightQ8_63_26_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_26_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_167 = _weightQ8_63_26_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_26_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_168 = _weightQ8_63_26_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_26_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_169 = _weightQ8_63_26_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_26_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_170 = _weightQ8_63_26_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_26_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_171 = _weightQ8_63_26_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_26_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_172 = _weightQ8_63_26_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_26_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_173 = _weightQ8_63_26_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_26_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_174 = _weightQ8_63_26_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_26_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_175 = _weightQ8_63_26_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_26_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_176 = _weightQ8_63_26_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_26_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_177 = _weightQ8_63_26_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_26_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_178 = _weightQ8_63_26_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_26_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_179 = _weightQ8_63_26_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_26_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_180 = _weightQ8_63_26_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_26_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_181 = _weightQ8_63_26_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_26_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_182 = _weightQ8_63_26_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_26_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_183 = _weightQ8_63_26_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_26_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_184 = _weightQ8_63_26_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_26_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_185 = _weightQ8_63_26_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_26_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_186 = _weightQ8_63_26_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_26_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_187 = _weightQ8_63_26_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_26_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_188 = _weightQ8_63_26_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_26_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_leadingZeros_T_189 = _weightQ8_63_26_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_26_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_26_leadingZeros = _weightQ8_63_26_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_26_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_26_expRaw_T_1 = 6'h1f - weightQ8_63_26_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_26_expRaw = weightQ8_63_26_isZero ? 6'h0 : _weightQ8_63_26_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_26_shiftAmt_T_2 = weightQ8_63_26_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_26_shiftAmt = weightQ8_63_26_expRaw > 6'h3 ? _weightQ8_63_26_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_26_mantissaRaw_T = weightQ8_63_26_absClipped >> weightQ8_63_26_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_26_mantissaRaw = _weightQ8_63_26_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_26_mantissa = weightQ8_63_26_expRaw >= 6'h3 ? weightQ8_63_26_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_26_expAdjusted = weightQ8_63_26_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_26_exp_T_4 = weightQ8_63_26_expAdjusted > 7'hf ? 4'hf : weightQ8_63_26_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_26_exp = weightQ8_63_26_isZero ? 4'h0 : _weightQ8_63_26_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_26_fp8 = {weightQ8_63_26_clippedX[31],weightQ8_63_26_exp,weightQ8_63_26_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_27_T = {24'h0,linear_weight_63_27}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_27_sign = _weightQ8_63_27_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_27_absX_T = ~_weightQ8_63_27_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_27_absX_T_2 = _weightQ8_63_27_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_27_absX = weightQ8_63_27_sign ? _weightQ8_63_27_absX_T_2 : _weightQ8_63_27_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_27_shiftedX_T_1 = _GEN_14432 - weightQ8_63_27_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_27_shiftedX_T_3 = weightQ8_63_27_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_27_shiftedX = weightQ8_63_27_sign ? _weightQ8_63_27_shiftedX_T_1 :
    _weightQ8_63_27_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_27_scaledX_T_1 = weightQ8_63_27_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_27_scaledX = _weightQ8_63_27_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_27_clippedX_T_2 = weightQ8_63_27_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_27_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_27_clippedX = weightQ8_63_27_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_27_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_27_absClipped_T_1 = ~weightQ8_63_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_27_absClipped_T_3 = _weightQ8_63_27_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_27_absClipped = weightQ8_63_27_clippedX[31] ? _weightQ8_63_27_absClipped_T_3 :
    weightQ8_63_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_27_isZero = weightQ8_63_27_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37611 = {{16'd0}, weightQ8_63_27_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_4 = _GEN_37611 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_6 = {weightQ8_63_27_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_8 = _weightQ8_63_27_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_9 = _weightQ8_63_27_leadingZeros_T_4 | _weightQ8_63_27_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37612 = {{8'd0}, _weightQ8_63_27_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_14 = _GEN_37612 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_16 = {_weightQ8_63_27_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_18 = _weightQ8_63_27_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_19 = _weightQ8_63_27_leadingZeros_T_14 | _weightQ8_63_27_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37613 = {{4'd0}, _weightQ8_63_27_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_24 = _GEN_37613 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_26 = {_weightQ8_63_27_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_28 = _weightQ8_63_27_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_29 = _weightQ8_63_27_leadingZeros_T_24 | _weightQ8_63_27_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37614 = {{2'd0}, _weightQ8_63_27_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_34 = _GEN_37614 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_36 = {_weightQ8_63_27_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_38 = _weightQ8_63_27_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_39 = _weightQ8_63_27_leadingZeros_T_34 | _weightQ8_63_27_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37615 = {{1'd0}, _weightQ8_63_27_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_44 = _GEN_37615 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_46 = {_weightQ8_63_27_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_48 = _weightQ8_63_27_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_27_leadingZeros_T_49 = _weightQ8_63_27_leadingZeros_T_44 | _weightQ8_63_27_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37616 = {{8'd0}, weightQ8_63_27_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_55 = _GEN_37616 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_57 = {weightQ8_63_27_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_59 = _weightQ8_63_27_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_60 = _weightQ8_63_27_leadingZeros_T_55 | _weightQ8_63_27_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37617 = {{4'd0}, _weightQ8_63_27_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_65 = _GEN_37617 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_67 = {_weightQ8_63_27_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_69 = _weightQ8_63_27_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_70 = _weightQ8_63_27_leadingZeros_T_65 | _weightQ8_63_27_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37618 = {{2'd0}, _weightQ8_63_27_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_75 = _GEN_37618 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_77 = {_weightQ8_63_27_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_79 = _weightQ8_63_27_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_80 = _weightQ8_63_27_leadingZeros_T_75 | _weightQ8_63_27_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37619 = {{1'd0}, _weightQ8_63_27_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_85 = _GEN_37619 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_87 = {_weightQ8_63_27_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_89 = _weightQ8_63_27_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_27_leadingZeros_T_90 = _weightQ8_63_27_leadingZeros_T_85 | _weightQ8_63_27_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_27_leadingZeros_T_93 = {_weightQ8_63_27_leadingZeros_T_49,_weightQ8_63_27_leadingZeros_T_90,
    weightQ8_63_27_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_143 = _weightQ8_63_27_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_144 = _weightQ8_63_27_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_27_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_145 = _weightQ8_63_27_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_27_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_146 = _weightQ8_63_27_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_27_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_147 = _weightQ8_63_27_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_27_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_148 = _weightQ8_63_27_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_27_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_149 = _weightQ8_63_27_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_27_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_150 = _weightQ8_63_27_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_27_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_151 = _weightQ8_63_27_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_27_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_152 = _weightQ8_63_27_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_27_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_153 = _weightQ8_63_27_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_27_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_154 = _weightQ8_63_27_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_27_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_155 = _weightQ8_63_27_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_27_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_156 = _weightQ8_63_27_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_27_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_157 = _weightQ8_63_27_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_27_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_158 = _weightQ8_63_27_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_27_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_159 = _weightQ8_63_27_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_27_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_160 = _weightQ8_63_27_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_27_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_161 = _weightQ8_63_27_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_27_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_162 = _weightQ8_63_27_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_27_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_163 = _weightQ8_63_27_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_27_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_164 = _weightQ8_63_27_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_27_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_165 = _weightQ8_63_27_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_27_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_166 = _weightQ8_63_27_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_27_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_167 = _weightQ8_63_27_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_27_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_168 = _weightQ8_63_27_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_27_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_169 = _weightQ8_63_27_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_27_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_170 = _weightQ8_63_27_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_27_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_171 = _weightQ8_63_27_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_27_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_172 = _weightQ8_63_27_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_27_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_173 = _weightQ8_63_27_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_27_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_174 = _weightQ8_63_27_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_27_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_175 = _weightQ8_63_27_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_27_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_176 = _weightQ8_63_27_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_27_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_177 = _weightQ8_63_27_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_27_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_178 = _weightQ8_63_27_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_27_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_179 = _weightQ8_63_27_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_27_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_180 = _weightQ8_63_27_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_27_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_181 = _weightQ8_63_27_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_27_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_182 = _weightQ8_63_27_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_27_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_183 = _weightQ8_63_27_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_27_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_184 = _weightQ8_63_27_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_27_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_185 = _weightQ8_63_27_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_27_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_186 = _weightQ8_63_27_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_27_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_187 = _weightQ8_63_27_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_27_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_188 = _weightQ8_63_27_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_27_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_leadingZeros_T_189 = _weightQ8_63_27_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_27_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_27_leadingZeros = _weightQ8_63_27_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_27_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_27_expRaw_T_1 = 6'h1f - weightQ8_63_27_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_27_expRaw = weightQ8_63_27_isZero ? 6'h0 : _weightQ8_63_27_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_27_shiftAmt_T_2 = weightQ8_63_27_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_27_shiftAmt = weightQ8_63_27_expRaw > 6'h3 ? _weightQ8_63_27_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_27_mantissaRaw_T = weightQ8_63_27_absClipped >> weightQ8_63_27_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_27_mantissaRaw = _weightQ8_63_27_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_27_mantissa = weightQ8_63_27_expRaw >= 6'h3 ? weightQ8_63_27_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_27_expAdjusted = weightQ8_63_27_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_27_exp_T_4 = weightQ8_63_27_expAdjusted > 7'hf ? 4'hf : weightQ8_63_27_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_27_exp = weightQ8_63_27_isZero ? 4'h0 : _weightQ8_63_27_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_27_fp8 = {weightQ8_63_27_clippedX[31],weightQ8_63_27_exp,weightQ8_63_27_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_28_T = {24'h0,linear_weight_63_28}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_28_sign = _weightQ8_63_28_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_28_absX_T = ~_weightQ8_63_28_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_28_absX_T_2 = _weightQ8_63_28_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_28_absX = weightQ8_63_28_sign ? _weightQ8_63_28_absX_T_2 : _weightQ8_63_28_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_28_shiftedX_T_1 = _GEN_14432 - weightQ8_63_28_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_28_shiftedX_T_3 = weightQ8_63_28_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_28_shiftedX = weightQ8_63_28_sign ? _weightQ8_63_28_shiftedX_T_1 :
    _weightQ8_63_28_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_28_scaledX_T_1 = weightQ8_63_28_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_28_scaledX = _weightQ8_63_28_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_28_clippedX_T_2 = weightQ8_63_28_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_28_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_28_clippedX = weightQ8_63_28_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_28_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_28_absClipped_T_1 = ~weightQ8_63_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_28_absClipped_T_3 = _weightQ8_63_28_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_28_absClipped = weightQ8_63_28_clippedX[31] ? _weightQ8_63_28_absClipped_T_3 :
    weightQ8_63_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_28_isZero = weightQ8_63_28_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37622 = {{16'd0}, weightQ8_63_28_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_4 = _GEN_37622 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_6 = {weightQ8_63_28_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_8 = _weightQ8_63_28_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_9 = _weightQ8_63_28_leadingZeros_T_4 | _weightQ8_63_28_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37623 = {{8'd0}, _weightQ8_63_28_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_14 = _GEN_37623 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_16 = {_weightQ8_63_28_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_18 = _weightQ8_63_28_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_19 = _weightQ8_63_28_leadingZeros_T_14 | _weightQ8_63_28_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37624 = {{4'd0}, _weightQ8_63_28_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_24 = _GEN_37624 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_26 = {_weightQ8_63_28_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_28 = _weightQ8_63_28_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_29 = _weightQ8_63_28_leadingZeros_T_24 | _weightQ8_63_28_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37625 = {{2'd0}, _weightQ8_63_28_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_34 = _GEN_37625 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_36 = {_weightQ8_63_28_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_38 = _weightQ8_63_28_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_39 = _weightQ8_63_28_leadingZeros_T_34 | _weightQ8_63_28_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37626 = {{1'd0}, _weightQ8_63_28_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_44 = _GEN_37626 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_46 = {_weightQ8_63_28_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_48 = _weightQ8_63_28_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_28_leadingZeros_T_49 = _weightQ8_63_28_leadingZeros_T_44 | _weightQ8_63_28_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37627 = {{8'd0}, weightQ8_63_28_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_55 = _GEN_37627 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_57 = {weightQ8_63_28_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_59 = _weightQ8_63_28_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_60 = _weightQ8_63_28_leadingZeros_T_55 | _weightQ8_63_28_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37628 = {{4'd0}, _weightQ8_63_28_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_65 = _GEN_37628 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_67 = {_weightQ8_63_28_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_69 = _weightQ8_63_28_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_70 = _weightQ8_63_28_leadingZeros_T_65 | _weightQ8_63_28_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37629 = {{2'd0}, _weightQ8_63_28_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_75 = _GEN_37629 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_77 = {_weightQ8_63_28_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_79 = _weightQ8_63_28_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_80 = _weightQ8_63_28_leadingZeros_T_75 | _weightQ8_63_28_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37630 = {{1'd0}, _weightQ8_63_28_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_85 = _GEN_37630 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_87 = {_weightQ8_63_28_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_89 = _weightQ8_63_28_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_28_leadingZeros_T_90 = _weightQ8_63_28_leadingZeros_T_85 | _weightQ8_63_28_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_28_leadingZeros_T_93 = {_weightQ8_63_28_leadingZeros_T_49,_weightQ8_63_28_leadingZeros_T_90,
    weightQ8_63_28_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_143 = _weightQ8_63_28_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_144 = _weightQ8_63_28_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_28_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_145 = _weightQ8_63_28_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_28_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_146 = _weightQ8_63_28_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_28_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_147 = _weightQ8_63_28_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_28_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_148 = _weightQ8_63_28_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_28_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_149 = _weightQ8_63_28_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_28_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_150 = _weightQ8_63_28_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_28_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_151 = _weightQ8_63_28_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_28_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_152 = _weightQ8_63_28_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_28_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_153 = _weightQ8_63_28_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_28_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_154 = _weightQ8_63_28_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_28_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_155 = _weightQ8_63_28_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_28_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_156 = _weightQ8_63_28_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_28_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_157 = _weightQ8_63_28_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_28_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_158 = _weightQ8_63_28_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_28_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_159 = _weightQ8_63_28_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_28_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_160 = _weightQ8_63_28_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_28_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_161 = _weightQ8_63_28_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_28_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_162 = _weightQ8_63_28_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_28_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_163 = _weightQ8_63_28_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_28_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_164 = _weightQ8_63_28_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_28_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_165 = _weightQ8_63_28_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_28_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_166 = _weightQ8_63_28_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_28_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_167 = _weightQ8_63_28_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_28_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_168 = _weightQ8_63_28_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_28_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_169 = _weightQ8_63_28_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_28_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_170 = _weightQ8_63_28_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_28_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_171 = _weightQ8_63_28_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_28_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_172 = _weightQ8_63_28_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_28_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_173 = _weightQ8_63_28_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_28_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_174 = _weightQ8_63_28_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_28_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_175 = _weightQ8_63_28_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_28_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_176 = _weightQ8_63_28_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_28_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_177 = _weightQ8_63_28_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_28_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_178 = _weightQ8_63_28_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_28_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_179 = _weightQ8_63_28_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_28_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_180 = _weightQ8_63_28_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_28_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_181 = _weightQ8_63_28_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_28_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_182 = _weightQ8_63_28_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_28_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_183 = _weightQ8_63_28_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_28_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_184 = _weightQ8_63_28_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_28_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_185 = _weightQ8_63_28_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_28_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_186 = _weightQ8_63_28_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_28_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_187 = _weightQ8_63_28_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_28_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_188 = _weightQ8_63_28_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_28_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_leadingZeros_T_189 = _weightQ8_63_28_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_28_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_28_leadingZeros = _weightQ8_63_28_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_28_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_28_expRaw_T_1 = 6'h1f - weightQ8_63_28_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_28_expRaw = weightQ8_63_28_isZero ? 6'h0 : _weightQ8_63_28_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_28_shiftAmt_T_2 = weightQ8_63_28_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_28_shiftAmt = weightQ8_63_28_expRaw > 6'h3 ? _weightQ8_63_28_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_28_mantissaRaw_T = weightQ8_63_28_absClipped >> weightQ8_63_28_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_28_mantissaRaw = _weightQ8_63_28_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_28_mantissa = weightQ8_63_28_expRaw >= 6'h3 ? weightQ8_63_28_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_28_expAdjusted = weightQ8_63_28_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_28_exp_T_4 = weightQ8_63_28_expAdjusted > 7'hf ? 4'hf : weightQ8_63_28_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_28_exp = weightQ8_63_28_isZero ? 4'h0 : _weightQ8_63_28_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_28_fp8 = {weightQ8_63_28_clippedX[31],weightQ8_63_28_exp,weightQ8_63_28_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_29_T = {24'h0,linear_weight_63_29}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_29_sign = _weightQ8_63_29_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_29_absX_T = ~_weightQ8_63_29_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_29_absX_T_2 = _weightQ8_63_29_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_29_absX = weightQ8_63_29_sign ? _weightQ8_63_29_absX_T_2 : _weightQ8_63_29_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_29_shiftedX_T_1 = _GEN_14432 - weightQ8_63_29_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_29_shiftedX_T_3 = weightQ8_63_29_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_29_shiftedX = weightQ8_63_29_sign ? _weightQ8_63_29_shiftedX_T_1 :
    _weightQ8_63_29_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_29_scaledX_T_1 = weightQ8_63_29_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_29_scaledX = _weightQ8_63_29_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_29_clippedX_T_2 = weightQ8_63_29_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_29_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_29_clippedX = weightQ8_63_29_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_29_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_29_absClipped_T_1 = ~weightQ8_63_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_29_absClipped_T_3 = _weightQ8_63_29_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_29_absClipped = weightQ8_63_29_clippedX[31] ? _weightQ8_63_29_absClipped_T_3 :
    weightQ8_63_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_29_isZero = weightQ8_63_29_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37633 = {{16'd0}, weightQ8_63_29_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_4 = _GEN_37633 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_6 = {weightQ8_63_29_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_8 = _weightQ8_63_29_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_9 = _weightQ8_63_29_leadingZeros_T_4 | _weightQ8_63_29_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37634 = {{8'd0}, _weightQ8_63_29_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_14 = _GEN_37634 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_16 = {_weightQ8_63_29_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_18 = _weightQ8_63_29_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_19 = _weightQ8_63_29_leadingZeros_T_14 | _weightQ8_63_29_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37635 = {{4'd0}, _weightQ8_63_29_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_24 = _GEN_37635 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_26 = {_weightQ8_63_29_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_28 = _weightQ8_63_29_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_29 = _weightQ8_63_29_leadingZeros_T_24 | _weightQ8_63_29_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37636 = {{2'd0}, _weightQ8_63_29_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_34 = _GEN_37636 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_36 = {_weightQ8_63_29_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_38 = _weightQ8_63_29_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_39 = _weightQ8_63_29_leadingZeros_T_34 | _weightQ8_63_29_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37637 = {{1'd0}, _weightQ8_63_29_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_44 = _GEN_37637 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_46 = {_weightQ8_63_29_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_48 = _weightQ8_63_29_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_29_leadingZeros_T_49 = _weightQ8_63_29_leadingZeros_T_44 | _weightQ8_63_29_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37638 = {{8'd0}, weightQ8_63_29_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_55 = _GEN_37638 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_57 = {weightQ8_63_29_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_59 = _weightQ8_63_29_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_60 = _weightQ8_63_29_leadingZeros_T_55 | _weightQ8_63_29_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37639 = {{4'd0}, _weightQ8_63_29_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_65 = _GEN_37639 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_67 = {_weightQ8_63_29_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_69 = _weightQ8_63_29_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_70 = _weightQ8_63_29_leadingZeros_T_65 | _weightQ8_63_29_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37640 = {{2'd0}, _weightQ8_63_29_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_75 = _GEN_37640 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_77 = {_weightQ8_63_29_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_79 = _weightQ8_63_29_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_80 = _weightQ8_63_29_leadingZeros_T_75 | _weightQ8_63_29_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37641 = {{1'd0}, _weightQ8_63_29_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_85 = _GEN_37641 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_87 = {_weightQ8_63_29_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_89 = _weightQ8_63_29_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_29_leadingZeros_T_90 = _weightQ8_63_29_leadingZeros_T_85 | _weightQ8_63_29_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_29_leadingZeros_T_93 = {_weightQ8_63_29_leadingZeros_T_49,_weightQ8_63_29_leadingZeros_T_90,
    weightQ8_63_29_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_143 = _weightQ8_63_29_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_144 = _weightQ8_63_29_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_29_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_145 = _weightQ8_63_29_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_29_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_146 = _weightQ8_63_29_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_29_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_147 = _weightQ8_63_29_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_29_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_148 = _weightQ8_63_29_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_29_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_149 = _weightQ8_63_29_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_29_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_150 = _weightQ8_63_29_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_29_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_151 = _weightQ8_63_29_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_29_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_152 = _weightQ8_63_29_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_29_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_153 = _weightQ8_63_29_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_29_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_154 = _weightQ8_63_29_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_29_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_155 = _weightQ8_63_29_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_29_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_156 = _weightQ8_63_29_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_29_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_157 = _weightQ8_63_29_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_29_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_158 = _weightQ8_63_29_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_29_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_159 = _weightQ8_63_29_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_29_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_160 = _weightQ8_63_29_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_29_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_161 = _weightQ8_63_29_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_29_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_162 = _weightQ8_63_29_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_29_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_163 = _weightQ8_63_29_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_29_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_164 = _weightQ8_63_29_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_29_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_165 = _weightQ8_63_29_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_29_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_166 = _weightQ8_63_29_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_29_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_167 = _weightQ8_63_29_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_29_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_168 = _weightQ8_63_29_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_29_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_169 = _weightQ8_63_29_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_29_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_170 = _weightQ8_63_29_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_29_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_171 = _weightQ8_63_29_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_29_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_172 = _weightQ8_63_29_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_29_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_173 = _weightQ8_63_29_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_29_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_174 = _weightQ8_63_29_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_29_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_175 = _weightQ8_63_29_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_29_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_176 = _weightQ8_63_29_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_29_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_177 = _weightQ8_63_29_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_29_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_178 = _weightQ8_63_29_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_29_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_179 = _weightQ8_63_29_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_29_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_180 = _weightQ8_63_29_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_29_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_181 = _weightQ8_63_29_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_29_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_182 = _weightQ8_63_29_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_29_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_183 = _weightQ8_63_29_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_29_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_184 = _weightQ8_63_29_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_29_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_185 = _weightQ8_63_29_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_29_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_186 = _weightQ8_63_29_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_29_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_187 = _weightQ8_63_29_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_29_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_188 = _weightQ8_63_29_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_29_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_leadingZeros_T_189 = _weightQ8_63_29_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_29_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_29_leadingZeros = _weightQ8_63_29_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_29_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_29_expRaw_T_1 = 6'h1f - weightQ8_63_29_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_29_expRaw = weightQ8_63_29_isZero ? 6'h0 : _weightQ8_63_29_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_29_shiftAmt_T_2 = weightQ8_63_29_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_29_shiftAmt = weightQ8_63_29_expRaw > 6'h3 ? _weightQ8_63_29_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_29_mantissaRaw_T = weightQ8_63_29_absClipped >> weightQ8_63_29_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_29_mantissaRaw = _weightQ8_63_29_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_29_mantissa = weightQ8_63_29_expRaw >= 6'h3 ? weightQ8_63_29_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_29_expAdjusted = weightQ8_63_29_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_29_exp_T_4 = weightQ8_63_29_expAdjusted > 7'hf ? 4'hf : weightQ8_63_29_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_29_exp = weightQ8_63_29_isZero ? 4'h0 : _weightQ8_63_29_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_29_fp8 = {weightQ8_63_29_clippedX[31],weightQ8_63_29_exp,weightQ8_63_29_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_30_T = {24'h0,linear_weight_63_30}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_30_sign = _weightQ8_63_30_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_30_absX_T = ~_weightQ8_63_30_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_30_absX_T_2 = _weightQ8_63_30_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_30_absX = weightQ8_63_30_sign ? _weightQ8_63_30_absX_T_2 : _weightQ8_63_30_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_30_shiftedX_T_1 = _GEN_14432 - weightQ8_63_30_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_30_shiftedX_T_3 = weightQ8_63_30_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_30_shiftedX = weightQ8_63_30_sign ? _weightQ8_63_30_shiftedX_T_1 :
    _weightQ8_63_30_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_30_scaledX_T_1 = weightQ8_63_30_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_30_scaledX = _weightQ8_63_30_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_30_clippedX_T_2 = weightQ8_63_30_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_30_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_30_clippedX = weightQ8_63_30_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_30_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_30_absClipped_T_1 = ~weightQ8_63_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_30_absClipped_T_3 = _weightQ8_63_30_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_30_absClipped = weightQ8_63_30_clippedX[31] ? _weightQ8_63_30_absClipped_T_3 :
    weightQ8_63_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_30_isZero = weightQ8_63_30_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37644 = {{16'd0}, weightQ8_63_30_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_4 = _GEN_37644 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_6 = {weightQ8_63_30_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_8 = _weightQ8_63_30_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_9 = _weightQ8_63_30_leadingZeros_T_4 | _weightQ8_63_30_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37645 = {{8'd0}, _weightQ8_63_30_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_14 = _GEN_37645 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_16 = {_weightQ8_63_30_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_18 = _weightQ8_63_30_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_19 = _weightQ8_63_30_leadingZeros_T_14 | _weightQ8_63_30_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37646 = {{4'd0}, _weightQ8_63_30_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_24 = _GEN_37646 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_26 = {_weightQ8_63_30_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_28 = _weightQ8_63_30_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_29 = _weightQ8_63_30_leadingZeros_T_24 | _weightQ8_63_30_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37647 = {{2'd0}, _weightQ8_63_30_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_34 = _GEN_37647 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_36 = {_weightQ8_63_30_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_38 = _weightQ8_63_30_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_39 = _weightQ8_63_30_leadingZeros_T_34 | _weightQ8_63_30_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37648 = {{1'd0}, _weightQ8_63_30_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_44 = _GEN_37648 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_46 = {_weightQ8_63_30_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_48 = _weightQ8_63_30_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_30_leadingZeros_T_49 = _weightQ8_63_30_leadingZeros_T_44 | _weightQ8_63_30_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37649 = {{8'd0}, weightQ8_63_30_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_55 = _GEN_37649 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_57 = {weightQ8_63_30_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_59 = _weightQ8_63_30_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_60 = _weightQ8_63_30_leadingZeros_T_55 | _weightQ8_63_30_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37650 = {{4'd0}, _weightQ8_63_30_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_65 = _GEN_37650 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_67 = {_weightQ8_63_30_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_69 = _weightQ8_63_30_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_70 = _weightQ8_63_30_leadingZeros_T_65 | _weightQ8_63_30_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37651 = {{2'd0}, _weightQ8_63_30_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_75 = _GEN_37651 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_77 = {_weightQ8_63_30_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_79 = _weightQ8_63_30_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_80 = _weightQ8_63_30_leadingZeros_T_75 | _weightQ8_63_30_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37652 = {{1'd0}, _weightQ8_63_30_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_85 = _GEN_37652 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_87 = {_weightQ8_63_30_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_89 = _weightQ8_63_30_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_30_leadingZeros_T_90 = _weightQ8_63_30_leadingZeros_T_85 | _weightQ8_63_30_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_30_leadingZeros_T_93 = {_weightQ8_63_30_leadingZeros_T_49,_weightQ8_63_30_leadingZeros_T_90,
    weightQ8_63_30_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_143 = _weightQ8_63_30_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_144 = _weightQ8_63_30_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_30_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_145 = _weightQ8_63_30_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_30_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_146 = _weightQ8_63_30_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_30_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_147 = _weightQ8_63_30_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_30_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_148 = _weightQ8_63_30_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_30_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_149 = _weightQ8_63_30_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_30_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_150 = _weightQ8_63_30_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_30_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_151 = _weightQ8_63_30_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_30_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_152 = _weightQ8_63_30_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_30_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_153 = _weightQ8_63_30_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_30_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_154 = _weightQ8_63_30_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_30_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_155 = _weightQ8_63_30_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_30_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_156 = _weightQ8_63_30_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_30_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_157 = _weightQ8_63_30_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_30_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_158 = _weightQ8_63_30_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_30_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_159 = _weightQ8_63_30_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_30_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_160 = _weightQ8_63_30_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_30_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_161 = _weightQ8_63_30_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_30_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_162 = _weightQ8_63_30_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_30_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_163 = _weightQ8_63_30_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_30_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_164 = _weightQ8_63_30_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_30_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_165 = _weightQ8_63_30_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_30_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_166 = _weightQ8_63_30_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_30_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_167 = _weightQ8_63_30_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_30_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_168 = _weightQ8_63_30_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_30_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_169 = _weightQ8_63_30_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_30_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_170 = _weightQ8_63_30_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_30_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_171 = _weightQ8_63_30_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_30_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_172 = _weightQ8_63_30_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_30_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_173 = _weightQ8_63_30_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_30_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_174 = _weightQ8_63_30_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_30_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_175 = _weightQ8_63_30_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_30_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_176 = _weightQ8_63_30_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_30_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_177 = _weightQ8_63_30_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_30_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_178 = _weightQ8_63_30_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_30_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_179 = _weightQ8_63_30_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_30_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_180 = _weightQ8_63_30_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_30_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_181 = _weightQ8_63_30_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_30_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_182 = _weightQ8_63_30_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_30_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_183 = _weightQ8_63_30_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_30_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_184 = _weightQ8_63_30_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_30_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_185 = _weightQ8_63_30_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_30_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_186 = _weightQ8_63_30_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_30_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_187 = _weightQ8_63_30_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_30_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_188 = _weightQ8_63_30_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_30_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_leadingZeros_T_189 = _weightQ8_63_30_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_30_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_30_leadingZeros = _weightQ8_63_30_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_30_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_30_expRaw_T_1 = 6'h1f - weightQ8_63_30_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_30_expRaw = weightQ8_63_30_isZero ? 6'h0 : _weightQ8_63_30_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_30_shiftAmt_T_2 = weightQ8_63_30_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_30_shiftAmt = weightQ8_63_30_expRaw > 6'h3 ? _weightQ8_63_30_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_30_mantissaRaw_T = weightQ8_63_30_absClipped >> weightQ8_63_30_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_30_mantissaRaw = _weightQ8_63_30_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_30_mantissa = weightQ8_63_30_expRaw >= 6'h3 ? weightQ8_63_30_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_30_expAdjusted = weightQ8_63_30_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_30_exp_T_4 = weightQ8_63_30_expAdjusted > 7'hf ? 4'hf : weightQ8_63_30_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_30_exp = weightQ8_63_30_isZero ? 4'h0 : _weightQ8_63_30_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_30_fp8 = {weightQ8_63_30_clippedX[31],weightQ8_63_30_exp,weightQ8_63_30_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] _weightQ8_63_31_T = {24'h0,linear_weight_63_31}; // @[src/main/scala/Multiple/LinearCompute.scala 118:49]
  wire  weightQ8_63_31_sign = _weightQ8_63_31_T[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _weightQ8_63_31_absX_T = ~_weightQ8_63_31_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _weightQ8_63_31_absX_T_2 = _weightQ8_63_31_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] weightQ8_63_31_absX = weightQ8_63_31_sign ? _weightQ8_63_31_absX_T_2 : _weightQ8_63_31_T; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _weightQ8_63_31_shiftedX_T_1 = _GEN_14432 - weightQ8_63_31_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _weightQ8_63_31_shiftedX_T_3 = weightQ8_63_31_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] weightQ8_63_31_shiftedX = weightQ8_63_31_sign ? _weightQ8_63_31_shiftedX_T_1 :
    _weightQ8_63_31_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _weightQ8_63_31_scaledX_T_1 = weightQ8_63_31_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] weightQ8_63_31_scaledX = _weightQ8_63_31_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _weightQ8_63_31_clippedX_T_2 = weightQ8_63_31_scaledX < 49'hfffffe40 ? 49'hfffffe40 :
    weightQ8_63_31_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] weightQ8_63_31_clippedX = weightQ8_63_31_scaledX > 49'h1c0 ? 49'h1c0 : _weightQ8_63_31_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _weightQ8_63_31_absClipped_T_1 = ~weightQ8_63_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _weightQ8_63_31_absClipped_T_3 = _weightQ8_63_31_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] weightQ8_63_31_absClipped = weightQ8_63_31_clippedX[31] ? _weightQ8_63_31_absClipped_T_3 :
    weightQ8_63_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  weightQ8_63_31_isZero = weightQ8_63_31_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_37655 = {{16'd0}, weightQ8_63_31_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_4 = _GEN_37655 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_6 = {weightQ8_63_31_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_8 = _weightQ8_63_31_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_9 = _weightQ8_63_31_leadingZeros_T_4 | _weightQ8_63_31_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37656 = {{8'd0}, _weightQ8_63_31_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_14 = _GEN_37656 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_16 = {_weightQ8_63_31_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_18 = _weightQ8_63_31_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_19 = _weightQ8_63_31_leadingZeros_T_14 | _weightQ8_63_31_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37657 = {{4'd0}, _weightQ8_63_31_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_24 = _GEN_37657 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_26 = {_weightQ8_63_31_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_28 = _weightQ8_63_31_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_29 = _weightQ8_63_31_leadingZeros_T_24 | _weightQ8_63_31_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37658 = {{2'd0}, _weightQ8_63_31_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_34 = _GEN_37658 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_36 = {_weightQ8_63_31_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_38 = _weightQ8_63_31_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_39 = _weightQ8_63_31_leadingZeros_T_34 | _weightQ8_63_31_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_37659 = {{1'd0}, _weightQ8_63_31_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_44 = _GEN_37659 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_46 = {_weightQ8_63_31_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_48 = _weightQ8_63_31_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _weightQ8_63_31_leadingZeros_T_49 = _weightQ8_63_31_leadingZeros_T_44 | _weightQ8_63_31_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37660 = {{8'd0}, weightQ8_63_31_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_55 = _GEN_37660 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_57 = {weightQ8_63_31_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_59 = _weightQ8_63_31_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_60 = _weightQ8_63_31_leadingZeros_T_55 | _weightQ8_63_31_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37661 = {{4'd0}, _weightQ8_63_31_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_65 = _GEN_37661 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_67 = {_weightQ8_63_31_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_69 = _weightQ8_63_31_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_70 = _weightQ8_63_31_leadingZeros_T_65 | _weightQ8_63_31_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37662 = {{2'd0}, _weightQ8_63_31_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_75 = _GEN_37662 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_77 = {_weightQ8_63_31_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_79 = _weightQ8_63_31_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_80 = _weightQ8_63_31_leadingZeros_T_75 | _weightQ8_63_31_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_37663 = {{1'd0}, _weightQ8_63_31_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_85 = _GEN_37663 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_87 = {_weightQ8_63_31_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_89 = _weightQ8_63_31_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _weightQ8_63_31_leadingZeros_T_90 = _weightQ8_63_31_leadingZeros_T_85 | _weightQ8_63_31_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _weightQ8_63_31_leadingZeros_T_93 = {_weightQ8_63_31_leadingZeros_T_49,_weightQ8_63_31_leadingZeros_T_90,
    weightQ8_63_31_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_143 = _weightQ8_63_31_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_144 = _weightQ8_63_31_leadingZeros_T_93[46] ? 6'h2e :
    _weightQ8_63_31_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_145 = _weightQ8_63_31_leadingZeros_T_93[45] ? 6'h2d :
    _weightQ8_63_31_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_146 = _weightQ8_63_31_leadingZeros_T_93[44] ? 6'h2c :
    _weightQ8_63_31_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_147 = _weightQ8_63_31_leadingZeros_T_93[43] ? 6'h2b :
    _weightQ8_63_31_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_148 = _weightQ8_63_31_leadingZeros_T_93[42] ? 6'h2a :
    _weightQ8_63_31_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_149 = _weightQ8_63_31_leadingZeros_T_93[41] ? 6'h29 :
    _weightQ8_63_31_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_150 = _weightQ8_63_31_leadingZeros_T_93[40] ? 6'h28 :
    _weightQ8_63_31_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_151 = _weightQ8_63_31_leadingZeros_T_93[39] ? 6'h27 :
    _weightQ8_63_31_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_152 = _weightQ8_63_31_leadingZeros_T_93[38] ? 6'h26 :
    _weightQ8_63_31_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_153 = _weightQ8_63_31_leadingZeros_T_93[37] ? 6'h25 :
    _weightQ8_63_31_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_154 = _weightQ8_63_31_leadingZeros_T_93[36] ? 6'h24 :
    _weightQ8_63_31_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_155 = _weightQ8_63_31_leadingZeros_T_93[35] ? 6'h23 :
    _weightQ8_63_31_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_156 = _weightQ8_63_31_leadingZeros_T_93[34] ? 6'h22 :
    _weightQ8_63_31_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_157 = _weightQ8_63_31_leadingZeros_T_93[33] ? 6'h21 :
    _weightQ8_63_31_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_158 = _weightQ8_63_31_leadingZeros_T_93[32] ? 6'h20 :
    _weightQ8_63_31_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_159 = _weightQ8_63_31_leadingZeros_T_93[31] ? 6'h1f :
    _weightQ8_63_31_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_160 = _weightQ8_63_31_leadingZeros_T_93[30] ? 6'h1e :
    _weightQ8_63_31_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_161 = _weightQ8_63_31_leadingZeros_T_93[29] ? 6'h1d :
    _weightQ8_63_31_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_162 = _weightQ8_63_31_leadingZeros_T_93[28] ? 6'h1c :
    _weightQ8_63_31_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_163 = _weightQ8_63_31_leadingZeros_T_93[27] ? 6'h1b :
    _weightQ8_63_31_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_164 = _weightQ8_63_31_leadingZeros_T_93[26] ? 6'h1a :
    _weightQ8_63_31_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_165 = _weightQ8_63_31_leadingZeros_T_93[25] ? 6'h19 :
    _weightQ8_63_31_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_166 = _weightQ8_63_31_leadingZeros_T_93[24] ? 6'h18 :
    _weightQ8_63_31_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_167 = _weightQ8_63_31_leadingZeros_T_93[23] ? 6'h17 :
    _weightQ8_63_31_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_168 = _weightQ8_63_31_leadingZeros_T_93[22] ? 6'h16 :
    _weightQ8_63_31_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_169 = _weightQ8_63_31_leadingZeros_T_93[21] ? 6'h15 :
    _weightQ8_63_31_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_170 = _weightQ8_63_31_leadingZeros_T_93[20] ? 6'h14 :
    _weightQ8_63_31_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_171 = _weightQ8_63_31_leadingZeros_T_93[19] ? 6'h13 :
    _weightQ8_63_31_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_172 = _weightQ8_63_31_leadingZeros_T_93[18] ? 6'h12 :
    _weightQ8_63_31_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_173 = _weightQ8_63_31_leadingZeros_T_93[17] ? 6'h11 :
    _weightQ8_63_31_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_174 = _weightQ8_63_31_leadingZeros_T_93[16] ? 6'h10 :
    _weightQ8_63_31_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_175 = _weightQ8_63_31_leadingZeros_T_93[15] ? 6'hf :
    _weightQ8_63_31_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_176 = _weightQ8_63_31_leadingZeros_T_93[14] ? 6'he :
    _weightQ8_63_31_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_177 = _weightQ8_63_31_leadingZeros_T_93[13] ? 6'hd :
    _weightQ8_63_31_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_178 = _weightQ8_63_31_leadingZeros_T_93[12] ? 6'hc :
    _weightQ8_63_31_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_179 = _weightQ8_63_31_leadingZeros_T_93[11] ? 6'hb :
    _weightQ8_63_31_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_180 = _weightQ8_63_31_leadingZeros_T_93[10] ? 6'ha :
    _weightQ8_63_31_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_181 = _weightQ8_63_31_leadingZeros_T_93[9] ? 6'h9 :
    _weightQ8_63_31_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_182 = _weightQ8_63_31_leadingZeros_T_93[8] ? 6'h8 :
    _weightQ8_63_31_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_183 = _weightQ8_63_31_leadingZeros_T_93[7] ? 6'h7 :
    _weightQ8_63_31_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_184 = _weightQ8_63_31_leadingZeros_T_93[6] ? 6'h6 :
    _weightQ8_63_31_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_185 = _weightQ8_63_31_leadingZeros_T_93[5] ? 6'h5 :
    _weightQ8_63_31_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_186 = _weightQ8_63_31_leadingZeros_T_93[4] ? 6'h4 :
    _weightQ8_63_31_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_187 = _weightQ8_63_31_leadingZeros_T_93[3] ? 6'h3 :
    _weightQ8_63_31_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_188 = _weightQ8_63_31_leadingZeros_T_93[2] ? 6'h2 :
    _weightQ8_63_31_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_leadingZeros_T_189 = _weightQ8_63_31_leadingZeros_T_93[1] ? 6'h1 :
    _weightQ8_63_31_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] weightQ8_63_31_leadingZeros = _weightQ8_63_31_leadingZeros_T_93[0] ? 6'h0 :
    _weightQ8_63_31_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _weightQ8_63_31_expRaw_T_1 = 6'h1f - weightQ8_63_31_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] weightQ8_63_31_expRaw = weightQ8_63_31_isZero ? 6'h0 : _weightQ8_63_31_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _weightQ8_63_31_shiftAmt_T_2 = weightQ8_63_31_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] weightQ8_63_31_shiftAmt = weightQ8_63_31_expRaw > 6'h3 ? _weightQ8_63_31_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _weightQ8_63_31_mantissaRaw_T = weightQ8_63_31_absClipped >> weightQ8_63_31_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] weightQ8_63_31_mantissaRaw = _weightQ8_63_31_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] weightQ8_63_31_mantissa = weightQ8_63_31_expRaw >= 6'h3 ? weightQ8_63_31_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] weightQ8_63_31_expAdjusted = weightQ8_63_31_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _weightQ8_63_31_exp_T_4 = weightQ8_63_31_expAdjusted > 7'hf ? 4'hf : weightQ8_63_31_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] weightQ8_63_31_exp = weightQ8_63_31_isZero ? 4'h0 : _weightQ8_63_31_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] weightQ8_63_31_fp8 = {weightQ8_63_31_clippedX[31],weightQ8_63_31_exp,weightQ8_63_31_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  reg [31:0] ansAll_63_0; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_1; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_2; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_3; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_4; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_5; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_6; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_7; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_8; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_9; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_10; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_11; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_12; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_13; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_14; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_15; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_16; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_17; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_18; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_19; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_20; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_21; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_22; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_23; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_24; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_25; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_26; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_27; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_28; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_29; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_30; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  reg [31:0] ansAll_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 123:21]
  wire  ansAll_63_0_signA = featuresInQ8_63[7]; // @[src/main/scala/Multiple/LinearCompute.scala 69:22]
  wire [3:0] ansAll_63_0_expA = featuresInQ8_63[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 70:21]
  wire [2:0] ansAll_63_0_mantA = featuresInQ8_63[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 71:22]
  wire  ansAll_63_0_signB = weightQ8_63_0[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_0_expB = weightQ8_63_0[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_0_mantB = weightQ8_63_0[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_0_mantissaA = {1'h1,ansAll_63_0_mantA}; // @[src/main/scala/Multiple/LinearCompute.scala 84:28]
  wire [3:0] ansAll_63_0_mantissaB = {1'h1,ansAll_63_0_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_0_expAUnbiased = ansAll_63_0_expA - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 87:33]
  wire [3:0] ansAll_63_0_expBUnbiased = ansAll_63_0_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_0_signProd = ansAll_63_0_signA ^ ansAll_63_0_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_0_mantProd = ansAll_63_0_mantissaA * ansAll_63_0_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_0_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_0_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_0_expProd = _ansAll_63_0_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_0_mantProdNorm = ansAll_63_0_mantProd[7] ? {{1'd0}, ansAll_63_0_mantProd[7:1]} :
    ansAll_63_0_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_0_expShift = {{3'd0}, ansAll_63_0_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39680 = {{1'd0}, ansAll_63_0_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_0_expFinal = ansAll_63_0_expProd + _GEN_39680; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_0 = {{31'd0}, ansAll_63_0_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_0_resultAbs_T_1 = _GEN_0 << ansAll_63_0_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_0_resultAbs = _ansAll_63_0_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_0_T_2 = ~ansAll_63_0_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_0_T_4 = _ansAll_63_0_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_1_signB = weightQ8_63_1[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_1_expB = weightQ8_63_1[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_1_mantB = weightQ8_63_1[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_1_mantissaB = {1'h1,ansAll_63_1_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_1_expBUnbiased = ansAll_63_1_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_1_signProd = ansAll_63_0_signA ^ ansAll_63_1_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_1_mantProd = ansAll_63_0_mantissaA * ansAll_63_1_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_1_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_1_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_1_expProd = _ansAll_63_1_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_1_mantProdNorm = ansAll_63_1_mantProd[7] ? {{1'd0}, ansAll_63_1_mantProd[7:1]} :
    ansAll_63_1_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_1_expShift = {{3'd0}, ansAll_63_1_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39681 = {{1'd0}, ansAll_63_1_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_1_expFinal = ansAll_63_1_expProd + _GEN_39681; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_1 = {{31'd0}, ansAll_63_1_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_1_resultAbs_T_1 = _GEN_1 << ansAll_63_1_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_1_resultAbs = _ansAll_63_1_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_1_T_2 = ~ansAll_63_1_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_1_T_4 = _ansAll_63_1_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_2_signB = weightQ8_63_2[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_2_expB = weightQ8_63_2[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_2_mantB = weightQ8_63_2[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_2_mantissaB = {1'h1,ansAll_63_2_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_2_expBUnbiased = ansAll_63_2_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_2_signProd = ansAll_63_0_signA ^ ansAll_63_2_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_2_mantProd = ansAll_63_0_mantissaA * ansAll_63_2_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_2_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_2_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_2_expProd = _ansAll_63_2_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_2_mantProdNorm = ansAll_63_2_mantProd[7] ? {{1'd0}, ansAll_63_2_mantProd[7:1]} :
    ansAll_63_2_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_2_expShift = {{3'd0}, ansAll_63_2_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39682 = {{1'd0}, ansAll_63_2_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_2_expFinal = ansAll_63_2_expProd + _GEN_39682; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_2 = {{31'd0}, ansAll_63_2_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_2_resultAbs_T_1 = _GEN_2 << ansAll_63_2_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_2_resultAbs = _ansAll_63_2_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_2_T_2 = ~ansAll_63_2_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_2_T_4 = _ansAll_63_2_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_3_signB = weightQ8_63_3[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_3_expB = weightQ8_63_3[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_3_mantB = weightQ8_63_3[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_3_mantissaB = {1'h1,ansAll_63_3_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_3_expBUnbiased = ansAll_63_3_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_3_signProd = ansAll_63_0_signA ^ ansAll_63_3_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_3_mantProd = ansAll_63_0_mantissaA * ansAll_63_3_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_3_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_3_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_3_expProd = _ansAll_63_3_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_3_mantProdNorm = ansAll_63_3_mantProd[7] ? {{1'd0}, ansAll_63_3_mantProd[7:1]} :
    ansAll_63_3_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_3_expShift = {{3'd0}, ansAll_63_3_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39683 = {{1'd0}, ansAll_63_3_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_3_expFinal = ansAll_63_3_expProd + _GEN_39683; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_3 = {{31'd0}, ansAll_63_3_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_3_resultAbs_T_1 = _GEN_3 << ansAll_63_3_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_3_resultAbs = _ansAll_63_3_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_3_T_2 = ~ansAll_63_3_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_3_T_4 = _ansAll_63_3_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_4_signB = weightQ8_63_4[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_4_expB = weightQ8_63_4[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_4_mantB = weightQ8_63_4[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_4_mantissaB = {1'h1,ansAll_63_4_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_4_expBUnbiased = ansAll_63_4_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_4_signProd = ansAll_63_0_signA ^ ansAll_63_4_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_4_mantProd = ansAll_63_0_mantissaA * ansAll_63_4_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_4_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_4_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_4_expProd = _ansAll_63_4_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_4_mantProdNorm = ansAll_63_4_mantProd[7] ? {{1'd0}, ansAll_63_4_mantProd[7:1]} :
    ansAll_63_4_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_4_expShift = {{3'd0}, ansAll_63_4_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39684 = {{1'd0}, ansAll_63_4_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_4_expFinal = ansAll_63_4_expProd + _GEN_39684; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_4 = {{31'd0}, ansAll_63_4_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_4_resultAbs_T_1 = _GEN_4 << ansAll_63_4_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_4_resultAbs = _ansAll_63_4_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_4_T_2 = ~ansAll_63_4_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_4_T_4 = _ansAll_63_4_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_5_signB = weightQ8_63_5[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_5_expB = weightQ8_63_5[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_5_mantB = weightQ8_63_5[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_5_mantissaB = {1'h1,ansAll_63_5_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_5_expBUnbiased = ansAll_63_5_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_5_signProd = ansAll_63_0_signA ^ ansAll_63_5_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_5_mantProd = ansAll_63_0_mantissaA * ansAll_63_5_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_5_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_5_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_5_expProd = _ansAll_63_5_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_5_mantProdNorm = ansAll_63_5_mantProd[7] ? {{1'd0}, ansAll_63_5_mantProd[7:1]} :
    ansAll_63_5_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_5_expShift = {{3'd0}, ansAll_63_5_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39685 = {{1'd0}, ansAll_63_5_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_5_expFinal = ansAll_63_5_expProd + _GEN_39685; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_5 = {{31'd0}, ansAll_63_5_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_5_resultAbs_T_1 = _GEN_5 << ansAll_63_5_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_5_resultAbs = _ansAll_63_5_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_5_T_2 = ~ansAll_63_5_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_5_T_4 = _ansAll_63_5_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_6_signB = weightQ8_63_6[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_6_expB = weightQ8_63_6[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_6_mantB = weightQ8_63_6[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_6_mantissaB = {1'h1,ansAll_63_6_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_6_expBUnbiased = ansAll_63_6_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_6_signProd = ansAll_63_0_signA ^ ansAll_63_6_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_6_mantProd = ansAll_63_0_mantissaA * ansAll_63_6_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_6_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_6_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_6_expProd = _ansAll_63_6_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_6_mantProdNorm = ansAll_63_6_mantProd[7] ? {{1'd0}, ansAll_63_6_mantProd[7:1]} :
    ansAll_63_6_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_6_expShift = {{3'd0}, ansAll_63_6_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39686 = {{1'd0}, ansAll_63_6_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_6_expFinal = ansAll_63_6_expProd + _GEN_39686; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_6 = {{31'd0}, ansAll_63_6_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_6_resultAbs_T_1 = _GEN_6 << ansAll_63_6_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_6_resultAbs = _ansAll_63_6_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_6_T_2 = ~ansAll_63_6_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_6_T_4 = _ansAll_63_6_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_7_signB = weightQ8_63_7[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_7_expB = weightQ8_63_7[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_7_mantB = weightQ8_63_7[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_7_mantissaB = {1'h1,ansAll_63_7_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_7_expBUnbiased = ansAll_63_7_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_7_signProd = ansAll_63_0_signA ^ ansAll_63_7_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_7_mantProd = ansAll_63_0_mantissaA * ansAll_63_7_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_7_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_7_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_7_expProd = _ansAll_63_7_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_7_mantProdNorm = ansAll_63_7_mantProd[7] ? {{1'd0}, ansAll_63_7_mantProd[7:1]} :
    ansAll_63_7_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_7_expShift = {{3'd0}, ansAll_63_7_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39687 = {{1'd0}, ansAll_63_7_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_7_expFinal = ansAll_63_7_expProd + _GEN_39687; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_7 = {{31'd0}, ansAll_63_7_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_7_resultAbs_T_1 = _GEN_7 << ansAll_63_7_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_7_resultAbs = _ansAll_63_7_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_7_T_2 = ~ansAll_63_7_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_7_T_4 = _ansAll_63_7_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_8_signB = weightQ8_63_8[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_8_expB = weightQ8_63_8[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_8_mantB = weightQ8_63_8[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_8_mantissaB = {1'h1,ansAll_63_8_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_8_expBUnbiased = ansAll_63_8_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_8_signProd = ansAll_63_0_signA ^ ansAll_63_8_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_8_mantProd = ansAll_63_0_mantissaA * ansAll_63_8_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_8_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_8_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_8_expProd = _ansAll_63_8_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_8_mantProdNorm = ansAll_63_8_mantProd[7] ? {{1'd0}, ansAll_63_8_mantProd[7:1]} :
    ansAll_63_8_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_8_expShift = {{3'd0}, ansAll_63_8_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39688 = {{1'd0}, ansAll_63_8_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_8_expFinal = ansAll_63_8_expProd + _GEN_39688; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_8 = {{31'd0}, ansAll_63_8_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_8_resultAbs_T_1 = _GEN_8 << ansAll_63_8_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_8_resultAbs = _ansAll_63_8_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_8_T_2 = ~ansAll_63_8_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_8_T_4 = _ansAll_63_8_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_9_signB = weightQ8_63_9[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_9_expB = weightQ8_63_9[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_9_mantB = weightQ8_63_9[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_9_mantissaB = {1'h1,ansAll_63_9_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_9_expBUnbiased = ansAll_63_9_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_9_signProd = ansAll_63_0_signA ^ ansAll_63_9_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_9_mantProd = ansAll_63_0_mantissaA * ansAll_63_9_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_9_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_9_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_9_expProd = _ansAll_63_9_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_9_mantProdNorm = ansAll_63_9_mantProd[7] ? {{1'd0}, ansAll_63_9_mantProd[7:1]} :
    ansAll_63_9_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_9_expShift = {{3'd0}, ansAll_63_9_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39689 = {{1'd0}, ansAll_63_9_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_9_expFinal = ansAll_63_9_expProd + _GEN_39689; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_9 = {{31'd0}, ansAll_63_9_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_9_resultAbs_T_1 = _GEN_9 << ansAll_63_9_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_9_resultAbs = _ansAll_63_9_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_9_T_2 = ~ansAll_63_9_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_9_T_4 = _ansAll_63_9_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_10_signB = weightQ8_63_10[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_10_expB = weightQ8_63_10[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_10_mantB = weightQ8_63_10[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_10_mantissaB = {1'h1,ansAll_63_10_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_10_expBUnbiased = ansAll_63_10_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_10_signProd = ansAll_63_0_signA ^ ansAll_63_10_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_10_mantProd = ansAll_63_0_mantissaA * ansAll_63_10_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_10_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_10_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_10_expProd = _ansAll_63_10_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_10_mantProdNorm = ansAll_63_10_mantProd[7] ? {{1'd0}, ansAll_63_10_mantProd[7:1]} :
    ansAll_63_10_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_10_expShift = {{3'd0}, ansAll_63_10_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39690 = {{1'd0}, ansAll_63_10_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_10_expFinal = ansAll_63_10_expProd + _GEN_39690; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_10 = {{31'd0}, ansAll_63_10_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_10_resultAbs_T_1 = _GEN_10 << ansAll_63_10_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_10_resultAbs = _ansAll_63_10_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_10_T_2 = ~ansAll_63_10_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_10_T_4 = _ansAll_63_10_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_11_signB = weightQ8_63_11[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_11_expB = weightQ8_63_11[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_11_mantB = weightQ8_63_11[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_11_mantissaB = {1'h1,ansAll_63_11_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_11_expBUnbiased = ansAll_63_11_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_11_signProd = ansAll_63_0_signA ^ ansAll_63_11_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_11_mantProd = ansAll_63_0_mantissaA * ansAll_63_11_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_11_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_11_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_11_expProd = _ansAll_63_11_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_11_mantProdNorm = ansAll_63_11_mantProd[7] ? {{1'd0}, ansAll_63_11_mantProd[7:1]} :
    ansAll_63_11_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_11_expShift = {{3'd0}, ansAll_63_11_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39691 = {{1'd0}, ansAll_63_11_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_11_expFinal = ansAll_63_11_expProd + _GEN_39691; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_11 = {{31'd0}, ansAll_63_11_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_11_resultAbs_T_1 = _GEN_11 << ansAll_63_11_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_11_resultAbs = _ansAll_63_11_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_11_T_2 = ~ansAll_63_11_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_11_T_4 = _ansAll_63_11_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_12_signB = weightQ8_63_12[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_12_expB = weightQ8_63_12[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_12_mantB = weightQ8_63_12[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_12_mantissaB = {1'h1,ansAll_63_12_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_12_expBUnbiased = ansAll_63_12_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_12_signProd = ansAll_63_0_signA ^ ansAll_63_12_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_12_mantProd = ansAll_63_0_mantissaA * ansAll_63_12_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_12_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_12_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_12_expProd = _ansAll_63_12_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_12_mantProdNorm = ansAll_63_12_mantProd[7] ? {{1'd0}, ansAll_63_12_mantProd[7:1]} :
    ansAll_63_12_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_12_expShift = {{3'd0}, ansAll_63_12_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39692 = {{1'd0}, ansAll_63_12_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_12_expFinal = ansAll_63_12_expProd + _GEN_39692; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_12 = {{31'd0}, ansAll_63_12_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_12_resultAbs_T_1 = _GEN_12 << ansAll_63_12_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_12_resultAbs = _ansAll_63_12_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_12_T_2 = ~ansAll_63_12_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_12_T_4 = _ansAll_63_12_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_13_signB = weightQ8_63_13[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_13_expB = weightQ8_63_13[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_13_mantB = weightQ8_63_13[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_13_mantissaB = {1'h1,ansAll_63_13_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_13_expBUnbiased = ansAll_63_13_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_13_signProd = ansAll_63_0_signA ^ ansAll_63_13_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_13_mantProd = ansAll_63_0_mantissaA * ansAll_63_13_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_13_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_13_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_13_expProd = _ansAll_63_13_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_13_mantProdNorm = ansAll_63_13_mantProd[7] ? {{1'd0}, ansAll_63_13_mantProd[7:1]} :
    ansAll_63_13_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_13_expShift = {{3'd0}, ansAll_63_13_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39693 = {{1'd0}, ansAll_63_13_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_13_expFinal = ansAll_63_13_expProd + _GEN_39693; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_13 = {{31'd0}, ansAll_63_13_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_13_resultAbs_T_1 = _GEN_13 << ansAll_63_13_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_13_resultAbs = _ansAll_63_13_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_13_T_2 = ~ansAll_63_13_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_13_T_4 = _ansAll_63_13_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_14_signB = weightQ8_63_14[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_14_expB = weightQ8_63_14[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_14_mantB = weightQ8_63_14[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_14_mantissaB = {1'h1,ansAll_63_14_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_14_expBUnbiased = ansAll_63_14_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_14_signProd = ansAll_63_0_signA ^ ansAll_63_14_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_14_mantProd = ansAll_63_0_mantissaA * ansAll_63_14_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_14_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_14_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_14_expProd = _ansAll_63_14_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_14_mantProdNorm = ansAll_63_14_mantProd[7] ? {{1'd0}, ansAll_63_14_mantProd[7:1]} :
    ansAll_63_14_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_14_expShift = {{3'd0}, ansAll_63_14_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39694 = {{1'd0}, ansAll_63_14_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_14_expFinal = ansAll_63_14_expProd + _GEN_39694; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_14 = {{31'd0}, ansAll_63_14_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_14_resultAbs_T_1 = _GEN_14 << ansAll_63_14_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_14_resultAbs = _ansAll_63_14_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_14_T_2 = ~ansAll_63_14_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_14_T_4 = _ansAll_63_14_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_15_signB = weightQ8_63_15[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_15_expB = weightQ8_63_15[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_15_mantB = weightQ8_63_15[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_15_mantissaB = {1'h1,ansAll_63_15_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_15_expBUnbiased = ansAll_63_15_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_15_signProd = ansAll_63_0_signA ^ ansAll_63_15_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_15_mantProd = ansAll_63_0_mantissaA * ansAll_63_15_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_15_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_15_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_15_expProd = _ansAll_63_15_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_15_mantProdNorm = ansAll_63_15_mantProd[7] ? {{1'd0}, ansAll_63_15_mantProd[7:1]} :
    ansAll_63_15_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_15_expShift = {{3'd0}, ansAll_63_15_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39695 = {{1'd0}, ansAll_63_15_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_15_expFinal = ansAll_63_15_expProd + _GEN_39695; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_15 = {{31'd0}, ansAll_63_15_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_15_resultAbs_T_1 = _GEN_15 << ansAll_63_15_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_15_resultAbs = _ansAll_63_15_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_15_T_2 = ~ansAll_63_15_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_15_T_4 = _ansAll_63_15_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_16_signB = weightQ8_63_16[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_16_expB = weightQ8_63_16[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_16_mantB = weightQ8_63_16[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_16_mantissaB = {1'h1,ansAll_63_16_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_16_expBUnbiased = ansAll_63_16_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_16_signProd = ansAll_63_0_signA ^ ansAll_63_16_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_16_mantProd = ansAll_63_0_mantissaA * ansAll_63_16_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_16_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_16_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_16_expProd = _ansAll_63_16_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_16_mantProdNorm = ansAll_63_16_mantProd[7] ? {{1'd0}, ansAll_63_16_mantProd[7:1]} :
    ansAll_63_16_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_16_expShift = {{3'd0}, ansAll_63_16_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39696 = {{1'd0}, ansAll_63_16_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_16_expFinal = ansAll_63_16_expProd + _GEN_39696; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_16 = {{31'd0}, ansAll_63_16_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_16_resultAbs_T_1 = _GEN_16 << ansAll_63_16_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_16_resultAbs = _ansAll_63_16_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_16_T_2 = ~ansAll_63_16_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_16_T_4 = _ansAll_63_16_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_17_signB = weightQ8_63_17[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_17_expB = weightQ8_63_17[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_17_mantB = weightQ8_63_17[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_17_mantissaB = {1'h1,ansAll_63_17_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_17_expBUnbiased = ansAll_63_17_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_17_signProd = ansAll_63_0_signA ^ ansAll_63_17_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_17_mantProd = ansAll_63_0_mantissaA * ansAll_63_17_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_17_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_17_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_17_expProd = _ansAll_63_17_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_17_mantProdNorm = ansAll_63_17_mantProd[7] ? {{1'd0}, ansAll_63_17_mantProd[7:1]} :
    ansAll_63_17_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_17_expShift = {{3'd0}, ansAll_63_17_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39697 = {{1'd0}, ansAll_63_17_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_17_expFinal = ansAll_63_17_expProd + _GEN_39697; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_17 = {{31'd0}, ansAll_63_17_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_17_resultAbs_T_1 = _GEN_17 << ansAll_63_17_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_17_resultAbs = _ansAll_63_17_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_17_T_2 = ~ansAll_63_17_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_17_T_4 = _ansAll_63_17_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_18_signB = weightQ8_63_18[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_18_expB = weightQ8_63_18[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_18_mantB = weightQ8_63_18[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_18_mantissaB = {1'h1,ansAll_63_18_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_18_expBUnbiased = ansAll_63_18_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_18_signProd = ansAll_63_0_signA ^ ansAll_63_18_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_18_mantProd = ansAll_63_0_mantissaA * ansAll_63_18_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_18_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_18_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_18_expProd = _ansAll_63_18_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_18_mantProdNorm = ansAll_63_18_mantProd[7] ? {{1'd0}, ansAll_63_18_mantProd[7:1]} :
    ansAll_63_18_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_18_expShift = {{3'd0}, ansAll_63_18_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39698 = {{1'd0}, ansAll_63_18_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_18_expFinal = ansAll_63_18_expProd + _GEN_39698; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_18 = {{31'd0}, ansAll_63_18_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_18_resultAbs_T_1 = _GEN_18 << ansAll_63_18_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_18_resultAbs = _ansAll_63_18_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_18_T_2 = ~ansAll_63_18_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_18_T_4 = _ansAll_63_18_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_19_signB = weightQ8_63_19[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_19_expB = weightQ8_63_19[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_19_mantB = weightQ8_63_19[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_19_mantissaB = {1'h1,ansAll_63_19_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_19_expBUnbiased = ansAll_63_19_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_19_signProd = ansAll_63_0_signA ^ ansAll_63_19_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_19_mantProd = ansAll_63_0_mantissaA * ansAll_63_19_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_19_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_19_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_19_expProd = _ansAll_63_19_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_19_mantProdNorm = ansAll_63_19_mantProd[7] ? {{1'd0}, ansAll_63_19_mantProd[7:1]} :
    ansAll_63_19_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_19_expShift = {{3'd0}, ansAll_63_19_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39699 = {{1'd0}, ansAll_63_19_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_19_expFinal = ansAll_63_19_expProd + _GEN_39699; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_19 = {{31'd0}, ansAll_63_19_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_19_resultAbs_T_1 = _GEN_19 << ansAll_63_19_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_19_resultAbs = _ansAll_63_19_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_19_T_2 = ~ansAll_63_19_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_19_T_4 = _ansAll_63_19_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_20_signB = weightQ8_63_20[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_20_expB = weightQ8_63_20[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_20_mantB = weightQ8_63_20[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_20_mantissaB = {1'h1,ansAll_63_20_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_20_expBUnbiased = ansAll_63_20_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_20_signProd = ansAll_63_0_signA ^ ansAll_63_20_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_20_mantProd = ansAll_63_0_mantissaA * ansAll_63_20_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_20_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_20_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_20_expProd = _ansAll_63_20_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_20_mantProdNorm = ansAll_63_20_mantProd[7] ? {{1'd0}, ansAll_63_20_mantProd[7:1]} :
    ansAll_63_20_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_20_expShift = {{3'd0}, ansAll_63_20_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39700 = {{1'd0}, ansAll_63_20_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_20_expFinal = ansAll_63_20_expProd + _GEN_39700; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_20 = {{31'd0}, ansAll_63_20_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_20_resultAbs_T_1 = _GEN_20 << ansAll_63_20_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_20_resultAbs = _ansAll_63_20_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_20_T_2 = ~ansAll_63_20_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_20_T_4 = _ansAll_63_20_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_21_signB = weightQ8_63_21[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_21_expB = weightQ8_63_21[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_21_mantB = weightQ8_63_21[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_21_mantissaB = {1'h1,ansAll_63_21_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_21_expBUnbiased = ansAll_63_21_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_21_signProd = ansAll_63_0_signA ^ ansAll_63_21_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_21_mantProd = ansAll_63_0_mantissaA * ansAll_63_21_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_21_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_21_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_21_expProd = _ansAll_63_21_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_21_mantProdNorm = ansAll_63_21_mantProd[7] ? {{1'd0}, ansAll_63_21_mantProd[7:1]} :
    ansAll_63_21_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_21_expShift = {{3'd0}, ansAll_63_21_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39701 = {{1'd0}, ansAll_63_21_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_21_expFinal = ansAll_63_21_expProd + _GEN_39701; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_21 = {{31'd0}, ansAll_63_21_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_21_resultAbs_T_1 = _GEN_21 << ansAll_63_21_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_21_resultAbs = _ansAll_63_21_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_21_T_2 = ~ansAll_63_21_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_21_T_4 = _ansAll_63_21_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_22_signB = weightQ8_63_22[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_22_expB = weightQ8_63_22[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_22_mantB = weightQ8_63_22[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_22_mantissaB = {1'h1,ansAll_63_22_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_22_expBUnbiased = ansAll_63_22_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_22_signProd = ansAll_63_0_signA ^ ansAll_63_22_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_22_mantProd = ansAll_63_0_mantissaA * ansAll_63_22_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_22_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_22_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_22_expProd = _ansAll_63_22_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_22_mantProdNorm = ansAll_63_22_mantProd[7] ? {{1'd0}, ansAll_63_22_mantProd[7:1]} :
    ansAll_63_22_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_22_expShift = {{3'd0}, ansAll_63_22_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39702 = {{1'd0}, ansAll_63_22_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_22_expFinal = ansAll_63_22_expProd + _GEN_39702; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_22 = {{31'd0}, ansAll_63_22_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_22_resultAbs_T_1 = _GEN_22 << ansAll_63_22_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_22_resultAbs = _ansAll_63_22_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_22_T_2 = ~ansAll_63_22_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_22_T_4 = _ansAll_63_22_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_23_signB = weightQ8_63_23[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_23_expB = weightQ8_63_23[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_23_mantB = weightQ8_63_23[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_23_mantissaB = {1'h1,ansAll_63_23_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_23_expBUnbiased = ansAll_63_23_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_23_signProd = ansAll_63_0_signA ^ ansAll_63_23_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_23_mantProd = ansAll_63_0_mantissaA * ansAll_63_23_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_23_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_23_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_23_expProd = _ansAll_63_23_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_23_mantProdNorm = ansAll_63_23_mantProd[7] ? {{1'd0}, ansAll_63_23_mantProd[7:1]} :
    ansAll_63_23_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_23_expShift = {{3'd0}, ansAll_63_23_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39703 = {{1'd0}, ansAll_63_23_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_23_expFinal = ansAll_63_23_expProd + _GEN_39703; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_23 = {{31'd0}, ansAll_63_23_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_23_resultAbs_T_1 = _GEN_23 << ansAll_63_23_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_23_resultAbs = _ansAll_63_23_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_23_T_2 = ~ansAll_63_23_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_23_T_4 = _ansAll_63_23_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_24_signB = weightQ8_63_24[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_24_expB = weightQ8_63_24[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_24_mantB = weightQ8_63_24[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_24_mantissaB = {1'h1,ansAll_63_24_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_24_expBUnbiased = ansAll_63_24_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_24_signProd = ansAll_63_0_signA ^ ansAll_63_24_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_24_mantProd = ansAll_63_0_mantissaA * ansAll_63_24_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_24_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_24_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_24_expProd = _ansAll_63_24_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_24_mantProdNorm = ansAll_63_24_mantProd[7] ? {{1'd0}, ansAll_63_24_mantProd[7:1]} :
    ansAll_63_24_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_24_expShift = {{3'd0}, ansAll_63_24_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39704 = {{1'd0}, ansAll_63_24_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_24_expFinal = ansAll_63_24_expProd + _GEN_39704; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_24 = {{31'd0}, ansAll_63_24_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_24_resultAbs_T_1 = _GEN_24 << ansAll_63_24_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_24_resultAbs = _ansAll_63_24_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_24_T_2 = ~ansAll_63_24_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_24_T_4 = _ansAll_63_24_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_25_signB = weightQ8_63_25[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_25_expB = weightQ8_63_25[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_25_mantB = weightQ8_63_25[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_25_mantissaB = {1'h1,ansAll_63_25_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_25_expBUnbiased = ansAll_63_25_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_25_signProd = ansAll_63_0_signA ^ ansAll_63_25_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_25_mantProd = ansAll_63_0_mantissaA * ansAll_63_25_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_25_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_25_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_25_expProd = _ansAll_63_25_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_25_mantProdNorm = ansAll_63_25_mantProd[7] ? {{1'd0}, ansAll_63_25_mantProd[7:1]} :
    ansAll_63_25_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_25_expShift = {{3'd0}, ansAll_63_25_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39705 = {{1'd0}, ansAll_63_25_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_25_expFinal = ansAll_63_25_expProd + _GEN_39705; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_25 = {{31'd0}, ansAll_63_25_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_25_resultAbs_T_1 = _GEN_25 << ansAll_63_25_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_25_resultAbs = _ansAll_63_25_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_25_T_2 = ~ansAll_63_25_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_25_T_4 = _ansAll_63_25_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_26_signB = weightQ8_63_26[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_26_expB = weightQ8_63_26[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_26_mantB = weightQ8_63_26[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_26_mantissaB = {1'h1,ansAll_63_26_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_26_expBUnbiased = ansAll_63_26_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_26_signProd = ansAll_63_0_signA ^ ansAll_63_26_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_26_mantProd = ansAll_63_0_mantissaA * ansAll_63_26_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_26_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_26_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_26_expProd = _ansAll_63_26_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_26_mantProdNorm = ansAll_63_26_mantProd[7] ? {{1'd0}, ansAll_63_26_mantProd[7:1]} :
    ansAll_63_26_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_26_expShift = {{3'd0}, ansAll_63_26_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39706 = {{1'd0}, ansAll_63_26_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_26_expFinal = ansAll_63_26_expProd + _GEN_39706; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_26 = {{31'd0}, ansAll_63_26_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_26_resultAbs_T_1 = _GEN_26 << ansAll_63_26_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_26_resultAbs = _ansAll_63_26_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_26_T_2 = ~ansAll_63_26_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_26_T_4 = _ansAll_63_26_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_27_signB = weightQ8_63_27[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_27_expB = weightQ8_63_27[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_27_mantB = weightQ8_63_27[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_27_mantissaB = {1'h1,ansAll_63_27_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_27_expBUnbiased = ansAll_63_27_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_27_signProd = ansAll_63_0_signA ^ ansAll_63_27_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_27_mantProd = ansAll_63_0_mantissaA * ansAll_63_27_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_27_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_27_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_27_expProd = _ansAll_63_27_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_27_mantProdNorm = ansAll_63_27_mantProd[7] ? {{1'd0}, ansAll_63_27_mantProd[7:1]} :
    ansAll_63_27_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_27_expShift = {{3'd0}, ansAll_63_27_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39707 = {{1'd0}, ansAll_63_27_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_27_expFinal = ansAll_63_27_expProd + _GEN_39707; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_27 = {{31'd0}, ansAll_63_27_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_27_resultAbs_T_1 = _GEN_27 << ansAll_63_27_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_27_resultAbs = _ansAll_63_27_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_27_T_2 = ~ansAll_63_27_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_27_T_4 = _ansAll_63_27_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_28_signB = weightQ8_63_28[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_28_expB = weightQ8_63_28[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_28_mantB = weightQ8_63_28[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_28_mantissaB = {1'h1,ansAll_63_28_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_28_expBUnbiased = ansAll_63_28_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_28_signProd = ansAll_63_0_signA ^ ansAll_63_28_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_28_mantProd = ansAll_63_0_mantissaA * ansAll_63_28_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_28_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_28_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_28_expProd = _ansAll_63_28_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_28_mantProdNorm = ansAll_63_28_mantProd[7] ? {{1'd0}, ansAll_63_28_mantProd[7:1]} :
    ansAll_63_28_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_28_expShift = {{3'd0}, ansAll_63_28_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39708 = {{1'd0}, ansAll_63_28_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_28_expFinal = ansAll_63_28_expProd + _GEN_39708; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_28 = {{31'd0}, ansAll_63_28_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_28_resultAbs_T_1 = _GEN_28 << ansAll_63_28_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_28_resultAbs = _ansAll_63_28_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_28_T_2 = ~ansAll_63_28_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_28_T_4 = _ansAll_63_28_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_29_signB = weightQ8_63_29[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_29_expB = weightQ8_63_29[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_29_mantB = weightQ8_63_29[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_29_mantissaB = {1'h1,ansAll_63_29_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_29_expBUnbiased = ansAll_63_29_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_29_signProd = ansAll_63_0_signA ^ ansAll_63_29_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_29_mantProd = ansAll_63_0_mantissaA * ansAll_63_29_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_29_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_29_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_29_expProd = _ansAll_63_29_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_29_mantProdNorm = ansAll_63_29_mantProd[7] ? {{1'd0}, ansAll_63_29_mantProd[7:1]} :
    ansAll_63_29_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_29_expShift = {{3'd0}, ansAll_63_29_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39709 = {{1'd0}, ansAll_63_29_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_29_expFinal = ansAll_63_29_expProd + _GEN_39709; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_29 = {{31'd0}, ansAll_63_29_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_29_resultAbs_T_1 = _GEN_29 << ansAll_63_29_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_29_resultAbs = _ansAll_63_29_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_29_T_2 = ~ansAll_63_29_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_29_T_4 = _ansAll_63_29_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_30_signB = weightQ8_63_30[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_30_expB = weightQ8_63_30[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_30_mantB = weightQ8_63_30[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_30_mantissaB = {1'h1,ansAll_63_30_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_30_expBUnbiased = ansAll_63_30_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_30_signProd = ansAll_63_0_signA ^ ansAll_63_30_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_30_mantProd = ansAll_63_0_mantissaA * ansAll_63_30_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_30_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_30_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_30_expProd = _ansAll_63_30_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_30_mantProdNorm = ansAll_63_30_mantProd[7] ? {{1'd0}, ansAll_63_30_mantProd[7:1]} :
    ansAll_63_30_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_30_expShift = {{3'd0}, ansAll_63_30_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39710 = {{1'd0}, ansAll_63_30_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_30_expFinal = ansAll_63_30_expProd + _GEN_39710; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_30 = {{31'd0}, ansAll_63_30_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_30_resultAbs_T_1 = _GEN_30 << ansAll_63_30_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_30_resultAbs = _ansAll_63_30_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_30_T_2 = ~ansAll_63_30_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_30_T_4 = _ansAll_63_30_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  wire  ansAll_63_31_signB = weightQ8_63_31[7]; // @[src/main/scala/Multiple/LinearCompute.scala 72:22]
  wire [3:0] ansAll_63_31_expB = weightQ8_63_31[6:3]; // @[src/main/scala/Multiple/LinearCompute.scala 73:21]
  wire [2:0] ansAll_63_31_mantB = weightQ8_63_31[2:0]; // @[src/main/scala/Multiple/LinearCompute.scala 74:22]
  wire [3:0] ansAll_63_31_mantissaB = {1'h1,ansAll_63_31_mantB}; // @[src/main/scala/Multiple/LinearCompute.scala 85:28]
  wire [3:0] ansAll_63_31_expBUnbiased = ansAll_63_31_expB - 4'h7; // @[src/main/scala/Multiple/LinearCompute.scala 88:33]
  wire  ansAll_63_31_signProd = ansAll_63_0_signA ^ ansAll_63_31_signB; // @[src/main/scala/Multiple/LinearCompute.scala 91:30]
  wire [7:0] ansAll_63_31_mantProd = ansAll_63_0_mantissaA * ansAll_63_31_mantissaB; // @[src/main/scala/Multiple/LinearCompute.scala 92:34]
  wire [4:0] _ansAll_63_31_expProd_T = ansAll_63_0_expAUnbiased + ansAll_63_31_expBUnbiased; // @[src/main/scala/Multiple/LinearCompute.scala 93:36]
  wire [4:0] ansAll_63_31_expProd = _ansAll_63_31_expProd_T + 5'h3; // @[src/main/scala/Multiple/LinearCompute.scala 93:52]
  wire [7:0] ansAll_63_31_mantProdNorm = ansAll_63_31_mantProd[7] ? {{1'd0}, ansAll_63_31_mantProd[7:1]} :
    ansAll_63_31_mantProd; // @[src/main/scala/Multiple/LinearCompute.scala 102:26 98:28 99:26]
  wire [3:0] ansAll_63_31_expShift = {{3'd0}, ansAll_63_31_mantProd[7]}; // @[src/main/scala/Multiple/LinearCompute.scala 97:28]
  wire [4:0] _GEN_39711 = {{1'd0}, ansAll_63_31_expShift}; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [4:0] ansAll_63_31_expFinal = ansAll_63_31_expProd + _GEN_39711; // @[src/main/scala/Multiple/LinearCompute.scala 106:32]
  wire [34:0] _GEN_31 = {{31'd0}, ansAll_63_31_mantProdNorm[6:3]}; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [34:0] _ansAll_63_31_resultAbs_T_1 = _GEN_31 << ansAll_63_31_expFinal; // @[src/main/scala/Multiple/LinearCompute.scala 107:45]
  wire [31:0] ansAll_63_31_resultAbs = _ansAll_63_31_resultAbs_T_1[31:0]; // @[src/main/scala/Multiple/LinearCompute.scala 107:57]
  wire [31:0] _ansAll_63_31_T_2 = ~ansAll_63_31_resultAbs; // @[src/main/scala/Multiple/LinearCompute.scala 110:24]
  wire [31:0] _ansAll_63_31_T_4 = _ansAll_63_31_T_2 + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 110:35]
  reg [7:0] ans_0; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_1; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_2; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_3; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_4; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_5; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_6; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_7; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_8; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_9; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_10; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_11; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_12; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_13; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_14; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_15; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_16; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_17; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_18; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_19; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_20; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_21; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_22; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_23; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_24; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_25; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_26; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_27; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_28; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_29; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_30; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [7:0] ans_31; // @[src/main/scala/Multiple/LinearCompute.scala 133:18]
  reg [31:0] tempSum_0; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_1; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_2; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_3; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_4; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_5; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_6; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_7; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_8; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_9; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_10; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_11; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_12; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_13; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_14; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_15; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_16; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_17; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_18; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_19; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_20; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_21; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_22; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_23; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_24; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_25; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_26; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_27; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_28; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_29; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_30; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  reg [31:0] tempSum_31; // @[src/main/scala/Multiple/LinearCompute.scala 134:22]
  wire [31:0] biasExtended = {24'h0,linear_bias_0}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32 = tempSum_0 + biasExtended; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_0_sign = sum32[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_0_absX_T = ~sum32; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_0_absX_T_2 = _ans_0_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_0_absX = ans_0_sign ? _ans_0_absX_T_2 : sum32; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_0_shiftedX_T_1 = _GEN_14432 - ans_0_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_0_shiftedX_T_3 = ans_0_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_0_shiftedX = ans_0_sign ? _ans_0_shiftedX_T_1 : _ans_0_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_0_scaledX_T_1 = ans_0_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_0_scaledX = _ans_0_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_0_clippedX_T_2 = ans_0_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_0_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_0_clippedX = ans_0_scaledX > 49'h1c0 ? 49'h1c0 : _ans_0_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_0_absClipped_T_1 = ~ans_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_0_absClipped_T_3 = _ans_0_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_0_absClipped = ans_0_clippedX[31] ? _ans_0_absClipped_T_3 : ans_0_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_0_isZero = ans_0_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39714 = {{16'd0}, ans_0_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_4 = _GEN_39714 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_6 = {ans_0_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_8 = _ans_0_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_9 = _ans_0_leadingZeros_T_4 | _ans_0_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39715 = {{8'd0}, _ans_0_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_14 = _GEN_39715 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_16 = {_ans_0_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_18 = _ans_0_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_19 = _ans_0_leadingZeros_T_14 | _ans_0_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39716 = {{4'd0}, _ans_0_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_24 = _GEN_39716 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_26 = {_ans_0_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_28 = _ans_0_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_29 = _ans_0_leadingZeros_T_24 | _ans_0_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39717 = {{2'd0}, _ans_0_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_34 = _GEN_39717 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_36 = {_ans_0_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_38 = _ans_0_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_39 = _ans_0_leadingZeros_T_34 | _ans_0_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39718 = {{1'd0}, _ans_0_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_44 = _GEN_39718 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_46 = {_ans_0_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_48 = _ans_0_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_0_leadingZeros_T_49 = _ans_0_leadingZeros_T_44 | _ans_0_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39719 = {{8'd0}, ans_0_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_55 = _GEN_39719 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_57 = {ans_0_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_59 = _ans_0_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_60 = _ans_0_leadingZeros_T_55 | _ans_0_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39720 = {{4'd0}, _ans_0_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_65 = _GEN_39720 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_67 = {_ans_0_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_69 = _ans_0_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_70 = _ans_0_leadingZeros_T_65 | _ans_0_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39721 = {{2'd0}, _ans_0_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_75 = _GEN_39721 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_77 = {_ans_0_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_79 = _ans_0_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_80 = _ans_0_leadingZeros_T_75 | _ans_0_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39722 = {{1'd0}, _ans_0_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_85 = _GEN_39722 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_87 = {_ans_0_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_89 = _ans_0_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_0_leadingZeros_T_90 = _ans_0_leadingZeros_T_85 | _ans_0_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_0_leadingZeros_T_93 = {_ans_0_leadingZeros_T_49,_ans_0_leadingZeros_T_90,ans_0_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_0_leadingZeros_T_143 = _ans_0_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_144 = _ans_0_leadingZeros_T_93[46] ? 6'h2e : _ans_0_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_145 = _ans_0_leadingZeros_T_93[45] ? 6'h2d : _ans_0_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_146 = _ans_0_leadingZeros_T_93[44] ? 6'h2c : _ans_0_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_147 = _ans_0_leadingZeros_T_93[43] ? 6'h2b : _ans_0_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_148 = _ans_0_leadingZeros_T_93[42] ? 6'h2a : _ans_0_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_149 = _ans_0_leadingZeros_T_93[41] ? 6'h29 : _ans_0_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_150 = _ans_0_leadingZeros_T_93[40] ? 6'h28 : _ans_0_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_151 = _ans_0_leadingZeros_T_93[39] ? 6'h27 : _ans_0_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_152 = _ans_0_leadingZeros_T_93[38] ? 6'h26 : _ans_0_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_153 = _ans_0_leadingZeros_T_93[37] ? 6'h25 : _ans_0_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_154 = _ans_0_leadingZeros_T_93[36] ? 6'h24 : _ans_0_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_155 = _ans_0_leadingZeros_T_93[35] ? 6'h23 : _ans_0_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_156 = _ans_0_leadingZeros_T_93[34] ? 6'h22 : _ans_0_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_157 = _ans_0_leadingZeros_T_93[33] ? 6'h21 : _ans_0_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_158 = _ans_0_leadingZeros_T_93[32] ? 6'h20 : _ans_0_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_159 = _ans_0_leadingZeros_T_93[31] ? 6'h1f : _ans_0_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_160 = _ans_0_leadingZeros_T_93[30] ? 6'h1e : _ans_0_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_161 = _ans_0_leadingZeros_T_93[29] ? 6'h1d : _ans_0_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_162 = _ans_0_leadingZeros_T_93[28] ? 6'h1c : _ans_0_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_163 = _ans_0_leadingZeros_T_93[27] ? 6'h1b : _ans_0_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_164 = _ans_0_leadingZeros_T_93[26] ? 6'h1a : _ans_0_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_165 = _ans_0_leadingZeros_T_93[25] ? 6'h19 : _ans_0_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_166 = _ans_0_leadingZeros_T_93[24] ? 6'h18 : _ans_0_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_167 = _ans_0_leadingZeros_T_93[23] ? 6'h17 : _ans_0_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_168 = _ans_0_leadingZeros_T_93[22] ? 6'h16 : _ans_0_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_169 = _ans_0_leadingZeros_T_93[21] ? 6'h15 : _ans_0_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_170 = _ans_0_leadingZeros_T_93[20] ? 6'h14 : _ans_0_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_171 = _ans_0_leadingZeros_T_93[19] ? 6'h13 : _ans_0_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_172 = _ans_0_leadingZeros_T_93[18] ? 6'h12 : _ans_0_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_173 = _ans_0_leadingZeros_T_93[17] ? 6'h11 : _ans_0_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_174 = _ans_0_leadingZeros_T_93[16] ? 6'h10 : _ans_0_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_175 = _ans_0_leadingZeros_T_93[15] ? 6'hf : _ans_0_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_176 = _ans_0_leadingZeros_T_93[14] ? 6'he : _ans_0_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_177 = _ans_0_leadingZeros_T_93[13] ? 6'hd : _ans_0_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_178 = _ans_0_leadingZeros_T_93[12] ? 6'hc : _ans_0_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_179 = _ans_0_leadingZeros_T_93[11] ? 6'hb : _ans_0_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_180 = _ans_0_leadingZeros_T_93[10] ? 6'ha : _ans_0_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_181 = _ans_0_leadingZeros_T_93[9] ? 6'h9 : _ans_0_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_182 = _ans_0_leadingZeros_T_93[8] ? 6'h8 : _ans_0_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_183 = _ans_0_leadingZeros_T_93[7] ? 6'h7 : _ans_0_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_184 = _ans_0_leadingZeros_T_93[6] ? 6'h6 : _ans_0_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_185 = _ans_0_leadingZeros_T_93[5] ? 6'h5 : _ans_0_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_186 = _ans_0_leadingZeros_T_93[4] ? 6'h4 : _ans_0_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_187 = _ans_0_leadingZeros_T_93[3] ? 6'h3 : _ans_0_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_188 = _ans_0_leadingZeros_T_93[2] ? 6'h2 : _ans_0_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_leadingZeros_T_189 = _ans_0_leadingZeros_T_93[1] ? 6'h1 : _ans_0_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_0_leadingZeros = _ans_0_leadingZeros_T_93[0] ? 6'h0 : _ans_0_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_0_expRaw_T_1 = 6'h1f - ans_0_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_0_expRaw = ans_0_isZero ? 6'h0 : _ans_0_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_0_shiftAmt_T_2 = ans_0_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_0_shiftAmt = ans_0_expRaw > 6'h3 ? _ans_0_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_0_mantissaRaw_T = ans_0_absClipped >> ans_0_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_0_mantissaRaw = _ans_0_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_0_mantissa = ans_0_expRaw >= 6'h3 ? ans_0_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_0_expAdjusted = ans_0_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_0_exp_T_4 = ans_0_expAdjusted > 7'hf ? 4'hf : ans_0_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_0_exp = ans_0_isZero ? 4'h0 : _ans_0_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_0_fp8 = {ans_0_clippedX[31],ans_0_exp,ans_0_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_1 = {24'h0,linear_bias_1}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_1 = tempSum_1 + biasExtended_1; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_1_sign = sum32_1[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_1_absX_T = ~sum32_1; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_1_absX_T_2 = _ans_1_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_1_absX = ans_1_sign ? _ans_1_absX_T_2 : sum32_1; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_1_shiftedX_T_1 = _GEN_14432 - ans_1_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_1_shiftedX_T_3 = ans_1_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_1_shiftedX = ans_1_sign ? _ans_1_shiftedX_T_1 : _ans_1_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_1_scaledX_T_1 = ans_1_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_1_scaledX = _ans_1_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_1_clippedX_T_2 = ans_1_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_1_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_1_clippedX = ans_1_scaledX > 49'h1c0 ? 49'h1c0 : _ans_1_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_1_absClipped_T_1 = ~ans_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_1_absClipped_T_3 = _ans_1_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_1_absClipped = ans_1_clippedX[31] ? _ans_1_absClipped_T_3 : ans_1_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_1_isZero = ans_1_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39725 = {{16'd0}, ans_1_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_4 = _GEN_39725 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_6 = {ans_1_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_8 = _ans_1_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_9 = _ans_1_leadingZeros_T_4 | _ans_1_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39726 = {{8'd0}, _ans_1_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_14 = _GEN_39726 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_16 = {_ans_1_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_18 = _ans_1_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_19 = _ans_1_leadingZeros_T_14 | _ans_1_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39727 = {{4'd0}, _ans_1_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_24 = _GEN_39727 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_26 = {_ans_1_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_28 = _ans_1_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_29 = _ans_1_leadingZeros_T_24 | _ans_1_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39728 = {{2'd0}, _ans_1_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_34 = _GEN_39728 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_36 = {_ans_1_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_38 = _ans_1_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_39 = _ans_1_leadingZeros_T_34 | _ans_1_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39729 = {{1'd0}, _ans_1_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_44 = _GEN_39729 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_46 = {_ans_1_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_48 = _ans_1_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_1_leadingZeros_T_49 = _ans_1_leadingZeros_T_44 | _ans_1_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39730 = {{8'd0}, ans_1_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_55 = _GEN_39730 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_57 = {ans_1_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_59 = _ans_1_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_60 = _ans_1_leadingZeros_T_55 | _ans_1_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39731 = {{4'd0}, _ans_1_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_65 = _GEN_39731 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_67 = {_ans_1_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_69 = _ans_1_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_70 = _ans_1_leadingZeros_T_65 | _ans_1_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39732 = {{2'd0}, _ans_1_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_75 = _GEN_39732 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_77 = {_ans_1_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_79 = _ans_1_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_80 = _ans_1_leadingZeros_T_75 | _ans_1_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39733 = {{1'd0}, _ans_1_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_85 = _GEN_39733 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_87 = {_ans_1_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_89 = _ans_1_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_1_leadingZeros_T_90 = _ans_1_leadingZeros_T_85 | _ans_1_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_1_leadingZeros_T_93 = {_ans_1_leadingZeros_T_49,_ans_1_leadingZeros_T_90,ans_1_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_1_leadingZeros_T_143 = _ans_1_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_144 = _ans_1_leadingZeros_T_93[46] ? 6'h2e : _ans_1_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_145 = _ans_1_leadingZeros_T_93[45] ? 6'h2d : _ans_1_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_146 = _ans_1_leadingZeros_T_93[44] ? 6'h2c : _ans_1_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_147 = _ans_1_leadingZeros_T_93[43] ? 6'h2b : _ans_1_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_148 = _ans_1_leadingZeros_T_93[42] ? 6'h2a : _ans_1_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_149 = _ans_1_leadingZeros_T_93[41] ? 6'h29 : _ans_1_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_150 = _ans_1_leadingZeros_T_93[40] ? 6'h28 : _ans_1_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_151 = _ans_1_leadingZeros_T_93[39] ? 6'h27 : _ans_1_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_152 = _ans_1_leadingZeros_T_93[38] ? 6'h26 : _ans_1_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_153 = _ans_1_leadingZeros_T_93[37] ? 6'h25 : _ans_1_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_154 = _ans_1_leadingZeros_T_93[36] ? 6'h24 : _ans_1_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_155 = _ans_1_leadingZeros_T_93[35] ? 6'h23 : _ans_1_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_156 = _ans_1_leadingZeros_T_93[34] ? 6'h22 : _ans_1_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_157 = _ans_1_leadingZeros_T_93[33] ? 6'h21 : _ans_1_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_158 = _ans_1_leadingZeros_T_93[32] ? 6'h20 : _ans_1_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_159 = _ans_1_leadingZeros_T_93[31] ? 6'h1f : _ans_1_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_160 = _ans_1_leadingZeros_T_93[30] ? 6'h1e : _ans_1_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_161 = _ans_1_leadingZeros_T_93[29] ? 6'h1d : _ans_1_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_162 = _ans_1_leadingZeros_T_93[28] ? 6'h1c : _ans_1_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_163 = _ans_1_leadingZeros_T_93[27] ? 6'h1b : _ans_1_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_164 = _ans_1_leadingZeros_T_93[26] ? 6'h1a : _ans_1_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_165 = _ans_1_leadingZeros_T_93[25] ? 6'h19 : _ans_1_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_166 = _ans_1_leadingZeros_T_93[24] ? 6'h18 : _ans_1_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_167 = _ans_1_leadingZeros_T_93[23] ? 6'h17 : _ans_1_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_168 = _ans_1_leadingZeros_T_93[22] ? 6'h16 : _ans_1_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_169 = _ans_1_leadingZeros_T_93[21] ? 6'h15 : _ans_1_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_170 = _ans_1_leadingZeros_T_93[20] ? 6'h14 : _ans_1_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_171 = _ans_1_leadingZeros_T_93[19] ? 6'h13 : _ans_1_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_172 = _ans_1_leadingZeros_T_93[18] ? 6'h12 : _ans_1_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_173 = _ans_1_leadingZeros_T_93[17] ? 6'h11 : _ans_1_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_174 = _ans_1_leadingZeros_T_93[16] ? 6'h10 : _ans_1_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_175 = _ans_1_leadingZeros_T_93[15] ? 6'hf : _ans_1_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_176 = _ans_1_leadingZeros_T_93[14] ? 6'he : _ans_1_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_177 = _ans_1_leadingZeros_T_93[13] ? 6'hd : _ans_1_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_178 = _ans_1_leadingZeros_T_93[12] ? 6'hc : _ans_1_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_179 = _ans_1_leadingZeros_T_93[11] ? 6'hb : _ans_1_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_180 = _ans_1_leadingZeros_T_93[10] ? 6'ha : _ans_1_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_181 = _ans_1_leadingZeros_T_93[9] ? 6'h9 : _ans_1_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_182 = _ans_1_leadingZeros_T_93[8] ? 6'h8 : _ans_1_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_183 = _ans_1_leadingZeros_T_93[7] ? 6'h7 : _ans_1_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_184 = _ans_1_leadingZeros_T_93[6] ? 6'h6 : _ans_1_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_185 = _ans_1_leadingZeros_T_93[5] ? 6'h5 : _ans_1_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_186 = _ans_1_leadingZeros_T_93[4] ? 6'h4 : _ans_1_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_187 = _ans_1_leadingZeros_T_93[3] ? 6'h3 : _ans_1_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_188 = _ans_1_leadingZeros_T_93[2] ? 6'h2 : _ans_1_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_leadingZeros_T_189 = _ans_1_leadingZeros_T_93[1] ? 6'h1 : _ans_1_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_1_leadingZeros = _ans_1_leadingZeros_T_93[0] ? 6'h0 : _ans_1_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_1_expRaw_T_1 = 6'h1f - ans_1_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_1_expRaw = ans_1_isZero ? 6'h0 : _ans_1_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_1_shiftAmt_T_2 = ans_1_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_1_shiftAmt = ans_1_expRaw > 6'h3 ? _ans_1_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_1_mantissaRaw_T = ans_1_absClipped >> ans_1_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_1_mantissaRaw = _ans_1_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_1_mantissa = ans_1_expRaw >= 6'h3 ? ans_1_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_1_expAdjusted = ans_1_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_1_exp_T_4 = ans_1_expAdjusted > 7'hf ? 4'hf : ans_1_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_1_exp = ans_1_isZero ? 4'h0 : _ans_1_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_1_fp8 = {ans_1_clippedX[31],ans_1_exp,ans_1_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_2 = {24'h0,linear_bias_2}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_2 = tempSum_2 + biasExtended_2; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_2_sign = sum32_2[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_2_absX_T = ~sum32_2; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_2_absX_T_2 = _ans_2_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_2_absX = ans_2_sign ? _ans_2_absX_T_2 : sum32_2; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_2_shiftedX_T_1 = _GEN_14432 - ans_2_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_2_shiftedX_T_3 = ans_2_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_2_shiftedX = ans_2_sign ? _ans_2_shiftedX_T_1 : _ans_2_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_2_scaledX_T_1 = ans_2_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_2_scaledX = _ans_2_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_2_clippedX_T_2 = ans_2_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_2_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_2_clippedX = ans_2_scaledX > 49'h1c0 ? 49'h1c0 : _ans_2_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_2_absClipped_T_1 = ~ans_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_2_absClipped_T_3 = _ans_2_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_2_absClipped = ans_2_clippedX[31] ? _ans_2_absClipped_T_3 : ans_2_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_2_isZero = ans_2_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39736 = {{16'd0}, ans_2_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_4 = _GEN_39736 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_6 = {ans_2_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_8 = _ans_2_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_9 = _ans_2_leadingZeros_T_4 | _ans_2_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39737 = {{8'd0}, _ans_2_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_14 = _GEN_39737 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_16 = {_ans_2_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_18 = _ans_2_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_19 = _ans_2_leadingZeros_T_14 | _ans_2_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39738 = {{4'd0}, _ans_2_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_24 = _GEN_39738 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_26 = {_ans_2_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_28 = _ans_2_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_29 = _ans_2_leadingZeros_T_24 | _ans_2_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39739 = {{2'd0}, _ans_2_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_34 = _GEN_39739 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_36 = {_ans_2_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_38 = _ans_2_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_39 = _ans_2_leadingZeros_T_34 | _ans_2_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39740 = {{1'd0}, _ans_2_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_44 = _GEN_39740 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_46 = {_ans_2_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_48 = _ans_2_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_2_leadingZeros_T_49 = _ans_2_leadingZeros_T_44 | _ans_2_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39741 = {{8'd0}, ans_2_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_55 = _GEN_39741 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_57 = {ans_2_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_59 = _ans_2_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_60 = _ans_2_leadingZeros_T_55 | _ans_2_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39742 = {{4'd0}, _ans_2_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_65 = _GEN_39742 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_67 = {_ans_2_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_69 = _ans_2_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_70 = _ans_2_leadingZeros_T_65 | _ans_2_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39743 = {{2'd0}, _ans_2_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_75 = _GEN_39743 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_77 = {_ans_2_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_79 = _ans_2_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_80 = _ans_2_leadingZeros_T_75 | _ans_2_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39744 = {{1'd0}, _ans_2_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_85 = _GEN_39744 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_87 = {_ans_2_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_89 = _ans_2_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_2_leadingZeros_T_90 = _ans_2_leadingZeros_T_85 | _ans_2_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_2_leadingZeros_T_93 = {_ans_2_leadingZeros_T_49,_ans_2_leadingZeros_T_90,ans_2_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_2_leadingZeros_T_143 = _ans_2_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_144 = _ans_2_leadingZeros_T_93[46] ? 6'h2e : _ans_2_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_145 = _ans_2_leadingZeros_T_93[45] ? 6'h2d : _ans_2_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_146 = _ans_2_leadingZeros_T_93[44] ? 6'h2c : _ans_2_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_147 = _ans_2_leadingZeros_T_93[43] ? 6'h2b : _ans_2_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_148 = _ans_2_leadingZeros_T_93[42] ? 6'h2a : _ans_2_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_149 = _ans_2_leadingZeros_T_93[41] ? 6'h29 : _ans_2_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_150 = _ans_2_leadingZeros_T_93[40] ? 6'h28 : _ans_2_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_151 = _ans_2_leadingZeros_T_93[39] ? 6'h27 : _ans_2_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_152 = _ans_2_leadingZeros_T_93[38] ? 6'h26 : _ans_2_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_153 = _ans_2_leadingZeros_T_93[37] ? 6'h25 : _ans_2_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_154 = _ans_2_leadingZeros_T_93[36] ? 6'h24 : _ans_2_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_155 = _ans_2_leadingZeros_T_93[35] ? 6'h23 : _ans_2_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_156 = _ans_2_leadingZeros_T_93[34] ? 6'h22 : _ans_2_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_157 = _ans_2_leadingZeros_T_93[33] ? 6'h21 : _ans_2_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_158 = _ans_2_leadingZeros_T_93[32] ? 6'h20 : _ans_2_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_159 = _ans_2_leadingZeros_T_93[31] ? 6'h1f : _ans_2_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_160 = _ans_2_leadingZeros_T_93[30] ? 6'h1e : _ans_2_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_161 = _ans_2_leadingZeros_T_93[29] ? 6'h1d : _ans_2_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_162 = _ans_2_leadingZeros_T_93[28] ? 6'h1c : _ans_2_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_163 = _ans_2_leadingZeros_T_93[27] ? 6'h1b : _ans_2_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_164 = _ans_2_leadingZeros_T_93[26] ? 6'h1a : _ans_2_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_165 = _ans_2_leadingZeros_T_93[25] ? 6'h19 : _ans_2_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_166 = _ans_2_leadingZeros_T_93[24] ? 6'h18 : _ans_2_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_167 = _ans_2_leadingZeros_T_93[23] ? 6'h17 : _ans_2_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_168 = _ans_2_leadingZeros_T_93[22] ? 6'h16 : _ans_2_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_169 = _ans_2_leadingZeros_T_93[21] ? 6'h15 : _ans_2_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_170 = _ans_2_leadingZeros_T_93[20] ? 6'h14 : _ans_2_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_171 = _ans_2_leadingZeros_T_93[19] ? 6'h13 : _ans_2_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_172 = _ans_2_leadingZeros_T_93[18] ? 6'h12 : _ans_2_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_173 = _ans_2_leadingZeros_T_93[17] ? 6'h11 : _ans_2_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_174 = _ans_2_leadingZeros_T_93[16] ? 6'h10 : _ans_2_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_175 = _ans_2_leadingZeros_T_93[15] ? 6'hf : _ans_2_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_176 = _ans_2_leadingZeros_T_93[14] ? 6'he : _ans_2_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_177 = _ans_2_leadingZeros_T_93[13] ? 6'hd : _ans_2_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_178 = _ans_2_leadingZeros_T_93[12] ? 6'hc : _ans_2_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_179 = _ans_2_leadingZeros_T_93[11] ? 6'hb : _ans_2_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_180 = _ans_2_leadingZeros_T_93[10] ? 6'ha : _ans_2_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_181 = _ans_2_leadingZeros_T_93[9] ? 6'h9 : _ans_2_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_182 = _ans_2_leadingZeros_T_93[8] ? 6'h8 : _ans_2_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_183 = _ans_2_leadingZeros_T_93[7] ? 6'h7 : _ans_2_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_184 = _ans_2_leadingZeros_T_93[6] ? 6'h6 : _ans_2_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_185 = _ans_2_leadingZeros_T_93[5] ? 6'h5 : _ans_2_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_186 = _ans_2_leadingZeros_T_93[4] ? 6'h4 : _ans_2_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_187 = _ans_2_leadingZeros_T_93[3] ? 6'h3 : _ans_2_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_188 = _ans_2_leadingZeros_T_93[2] ? 6'h2 : _ans_2_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_leadingZeros_T_189 = _ans_2_leadingZeros_T_93[1] ? 6'h1 : _ans_2_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_2_leadingZeros = _ans_2_leadingZeros_T_93[0] ? 6'h0 : _ans_2_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_2_expRaw_T_1 = 6'h1f - ans_2_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_2_expRaw = ans_2_isZero ? 6'h0 : _ans_2_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_2_shiftAmt_T_2 = ans_2_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_2_shiftAmt = ans_2_expRaw > 6'h3 ? _ans_2_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_2_mantissaRaw_T = ans_2_absClipped >> ans_2_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_2_mantissaRaw = _ans_2_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_2_mantissa = ans_2_expRaw >= 6'h3 ? ans_2_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_2_expAdjusted = ans_2_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_2_exp_T_4 = ans_2_expAdjusted > 7'hf ? 4'hf : ans_2_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_2_exp = ans_2_isZero ? 4'h0 : _ans_2_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_2_fp8 = {ans_2_clippedX[31],ans_2_exp,ans_2_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_3 = {24'h0,linear_bias_3}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_3 = tempSum_3 + biasExtended_3; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_3_sign = sum32_3[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_3_absX_T = ~sum32_3; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_3_absX_T_2 = _ans_3_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_3_absX = ans_3_sign ? _ans_3_absX_T_2 : sum32_3; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_3_shiftedX_T_1 = _GEN_14432 - ans_3_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_3_shiftedX_T_3 = ans_3_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_3_shiftedX = ans_3_sign ? _ans_3_shiftedX_T_1 : _ans_3_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_3_scaledX_T_1 = ans_3_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_3_scaledX = _ans_3_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_3_clippedX_T_2 = ans_3_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_3_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_3_clippedX = ans_3_scaledX > 49'h1c0 ? 49'h1c0 : _ans_3_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_3_absClipped_T_1 = ~ans_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_3_absClipped_T_3 = _ans_3_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_3_absClipped = ans_3_clippedX[31] ? _ans_3_absClipped_T_3 : ans_3_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_3_isZero = ans_3_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39747 = {{16'd0}, ans_3_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_4 = _GEN_39747 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_6 = {ans_3_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_8 = _ans_3_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_9 = _ans_3_leadingZeros_T_4 | _ans_3_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39748 = {{8'd0}, _ans_3_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_14 = _GEN_39748 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_16 = {_ans_3_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_18 = _ans_3_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_19 = _ans_3_leadingZeros_T_14 | _ans_3_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39749 = {{4'd0}, _ans_3_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_24 = _GEN_39749 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_26 = {_ans_3_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_28 = _ans_3_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_29 = _ans_3_leadingZeros_T_24 | _ans_3_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39750 = {{2'd0}, _ans_3_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_34 = _GEN_39750 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_36 = {_ans_3_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_38 = _ans_3_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_39 = _ans_3_leadingZeros_T_34 | _ans_3_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39751 = {{1'd0}, _ans_3_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_44 = _GEN_39751 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_46 = {_ans_3_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_48 = _ans_3_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_3_leadingZeros_T_49 = _ans_3_leadingZeros_T_44 | _ans_3_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39752 = {{8'd0}, ans_3_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_55 = _GEN_39752 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_57 = {ans_3_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_59 = _ans_3_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_60 = _ans_3_leadingZeros_T_55 | _ans_3_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39753 = {{4'd0}, _ans_3_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_65 = _GEN_39753 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_67 = {_ans_3_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_69 = _ans_3_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_70 = _ans_3_leadingZeros_T_65 | _ans_3_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39754 = {{2'd0}, _ans_3_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_75 = _GEN_39754 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_77 = {_ans_3_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_79 = _ans_3_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_80 = _ans_3_leadingZeros_T_75 | _ans_3_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39755 = {{1'd0}, _ans_3_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_85 = _GEN_39755 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_87 = {_ans_3_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_89 = _ans_3_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_3_leadingZeros_T_90 = _ans_3_leadingZeros_T_85 | _ans_3_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_3_leadingZeros_T_93 = {_ans_3_leadingZeros_T_49,_ans_3_leadingZeros_T_90,ans_3_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_3_leadingZeros_T_143 = _ans_3_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_144 = _ans_3_leadingZeros_T_93[46] ? 6'h2e : _ans_3_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_145 = _ans_3_leadingZeros_T_93[45] ? 6'h2d : _ans_3_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_146 = _ans_3_leadingZeros_T_93[44] ? 6'h2c : _ans_3_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_147 = _ans_3_leadingZeros_T_93[43] ? 6'h2b : _ans_3_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_148 = _ans_3_leadingZeros_T_93[42] ? 6'h2a : _ans_3_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_149 = _ans_3_leadingZeros_T_93[41] ? 6'h29 : _ans_3_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_150 = _ans_3_leadingZeros_T_93[40] ? 6'h28 : _ans_3_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_151 = _ans_3_leadingZeros_T_93[39] ? 6'h27 : _ans_3_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_152 = _ans_3_leadingZeros_T_93[38] ? 6'h26 : _ans_3_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_153 = _ans_3_leadingZeros_T_93[37] ? 6'h25 : _ans_3_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_154 = _ans_3_leadingZeros_T_93[36] ? 6'h24 : _ans_3_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_155 = _ans_3_leadingZeros_T_93[35] ? 6'h23 : _ans_3_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_156 = _ans_3_leadingZeros_T_93[34] ? 6'h22 : _ans_3_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_157 = _ans_3_leadingZeros_T_93[33] ? 6'h21 : _ans_3_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_158 = _ans_3_leadingZeros_T_93[32] ? 6'h20 : _ans_3_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_159 = _ans_3_leadingZeros_T_93[31] ? 6'h1f : _ans_3_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_160 = _ans_3_leadingZeros_T_93[30] ? 6'h1e : _ans_3_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_161 = _ans_3_leadingZeros_T_93[29] ? 6'h1d : _ans_3_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_162 = _ans_3_leadingZeros_T_93[28] ? 6'h1c : _ans_3_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_163 = _ans_3_leadingZeros_T_93[27] ? 6'h1b : _ans_3_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_164 = _ans_3_leadingZeros_T_93[26] ? 6'h1a : _ans_3_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_165 = _ans_3_leadingZeros_T_93[25] ? 6'h19 : _ans_3_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_166 = _ans_3_leadingZeros_T_93[24] ? 6'h18 : _ans_3_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_167 = _ans_3_leadingZeros_T_93[23] ? 6'h17 : _ans_3_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_168 = _ans_3_leadingZeros_T_93[22] ? 6'h16 : _ans_3_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_169 = _ans_3_leadingZeros_T_93[21] ? 6'h15 : _ans_3_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_170 = _ans_3_leadingZeros_T_93[20] ? 6'h14 : _ans_3_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_171 = _ans_3_leadingZeros_T_93[19] ? 6'h13 : _ans_3_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_172 = _ans_3_leadingZeros_T_93[18] ? 6'h12 : _ans_3_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_173 = _ans_3_leadingZeros_T_93[17] ? 6'h11 : _ans_3_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_174 = _ans_3_leadingZeros_T_93[16] ? 6'h10 : _ans_3_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_175 = _ans_3_leadingZeros_T_93[15] ? 6'hf : _ans_3_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_176 = _ans_3_leadingZeros_T_93[14] ? 6'he : _ans_3_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_177 = _ans_3_leadingZeros_T_93[13] ? 6'hd : _ans_3_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_178 = _ans_3_leadingZeros_T_93[12] ? 6'hc : _ans_3_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_179 = _ans_3_leadingZeros_T_93[11] ? 6'hb : _ans_3_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_180 = _ans_3_leadingZeros_T_93[10] ? 6'ha : _ans_3_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_181 = _ans_3_leadingZeros_T_93[9] ? 6'h9 : _ans_3_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_182 = _ans_3_leadingZeros_T_93[8] ? 6'h8 : _ans_3_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_183 = _ans_3_leadingZeros_T_93[7] ? 6'h7 : _ans_3_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_184 = _ans_3_leadingZeros_T_93[6] ? 6'h6 : _ans_3_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_185 = _ans_3_leadingZeros_T_93[5] ? 6'h5 : _ans_3_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_186 = _ans_3_leadingZeros_T_93[4] ? 6'h4 : _ans_3_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_187 = _ans_3_leadingZeros_T_93[3] ? 6'h3 : _ans_3_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_188 = _ans_3_leadingZeros_T_93[2] ? 6'h2 : _ans_3_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_leadingZeros_T_189 = _ans_3_leadingZeros_T_93[1] ? 6'h1 : _ans_3_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_3_leadingZeros = _ans_3_leadingZeros_T_93[0] ? 6'h0 : _ans_3_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_3_expRaw_T_1 = 6'h1f - ans_3_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_3_expRaw = ans_3_isZero ? 6'h0 : _ans_3_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_3_shiftAmt_T_2 = ans_3_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_3_shiftAmt = ans_3_expRaw > 6'h3 ? _ans_3_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_3_mantissaRaw_T = ans_3_absClipped >> ans_3_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_3_mantissaRaw = _ans_3_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_3_mantissa = ans_3_expRaw >= 6'h3 ? ans_3_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_3_expAdjusted = ans_3_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_3_exp_T_4 = ans_3_expAdjusted > 7'hf ? 4'hf : ans_3_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_3_exp = ans_3_isZero ? 4'h0 : _ans_3_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_3_fp8 = {ans_3_clippedX[31],ans_3_exp,ans_3_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_4 = {24'h0,linear_bias_4}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_4 = tempSum_4 + biasExtended_4; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_4_sign = sum32_4[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_4_absX_T = ~sum32_4; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_4_absX_T_2 = _ans_4_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_4_absX = ans_4_sign ? _ans_4_absX_T_2 : sum32_4; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_4_shiftedX_T_1 = _GEN_14432 - ans_4_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_4_shiftedX_T_3 = ans_4_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_4_shiftedX = ans_4_sign ? _ans_4_shiftedX_T_1 : _ans_4_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_4_scaledX_T_1 = ans_4_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_4_scaledX = _ans_4_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_4_clippedX_T_2 = ans_4_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_4_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_4_clippedX = ans_4_scaledX > 49'h1c0 ? 49'h1c0 : _ans_4_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_4_absClipped_T_1 = ~ans_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_4_absClipped_T_3 = _ans_4_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_4_absClipped = ans_4_clippedX[31] ? _ans_4_absClipped_T_3 : ans_4_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_4_isZero = ans_4_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39758 = {{16'd0}, ans_4_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_4 = _GEN_39758 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_6 = {ans_4_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_8 = _ans_4_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_9 = _ans_4_leadingZeros_T_4 | _ans_4_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39759 = {{8'd0}, _ans_4_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_14 = _GEN_39759 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_16 = {_ans_4_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_18 = _ans_4_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_19 = _ans_4_leadingZeros_T_14 | _ans_4_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39760 = {{4'd0}, _ans_4_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_24 = _GEN_39760 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_26 = {_ans_4_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_28 = _ans_4_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_29 = _ans_4_leadingZeros_T_24 | _ans_4_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39761 = {{2'd0}, _ans_4_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_34 = _GEN_39761 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_36 = {_ans_4_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_38 = _ans_4_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_39 = _ans_4_leadingZeros_T_34 | _ans_4_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39762 = {{1'd0}, _ans_4_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_44 = _GEN_39762 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_46 = {_ans_4_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_48 = _ans_4_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_4_leadingZeros_T_49 = _ans_4_leadingZeros_T_44 | _ans_4_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39763 = {{8'd0}, ans_4_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_55 = _GEN_39763 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_57 = {ans_4_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_59 = _ans_4_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_60 = _ans_4_leadingZeros_T_55 | _ans_4_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39764 = {{4'd0}, _ans_4_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_65 = _GEN_39764 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_67 = {_ans_4_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_69 = _ans_4_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_70 = _ans_4_leadingZeros_T_65 | _ans_4_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39765 = {{2'd0}, _ans_4_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_75 = _GEN_39765 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_77 = {_ans_4_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_79 = _ans_4_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_80 = _ans_4_leadingZeros_T_75 | _ans_4_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39766 = {{1'd0}, _ans_4_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_85 = _GEN_39766 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_87 = {_ans_4_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_89 = _ans_4_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_4_leadingZeros_T_90 = _ans_4_leadingZeros_T_85 | _ans_4_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_4_leadingZeros_T_93 = {_ans_4_leadingZeros_T_49,_ans_4_leadingZeros_T_90,ans_4_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_4_leadingZeros_T_143 = _ans_4_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_144 = _ans_4_leadingZeros_T_93[46] ? 6'h2e : _ans_4_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_145 = _ans_4_leadingZeros_T_93[45] ? 6'h2d : _ans_4_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_146 = _ans_4_leadingZeros_T_93[44] ? 6'h2c : _ans_4_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_147 = _ans_4_leadingZeros_T_93[43] ? 6'h2b : _ans_4_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_148 = _ans_4_leadingZeros_T_93[42] ? 6'h2a : _ans_4_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_149 = _ans_4_leadingZeros_T_93[41] ? 6'h29 : _ans_4_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_150 = _ans_4_leadingZeros_T_93[40] ? 6'h28 : _ans_4_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_151 = _ans_4_leadingZeros_T_93[39] ? 6'h27 : _ans_4_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_152 = _ans_4_leadingZeros_T_93[38] ? 6'h26 : _ans_4_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_153 = _ans_4_leadingZeros_T_93[37] ? 6'h25 : _ans_4_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_154 = _ans_4_leadingZeros_T_93[36] ? 6'h24 : _ans_4_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_155 = _ans_4_leadingZeros_T_93[35] ? 6'h23 : _ans_4_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_156 = _ans_4_leadingZeros_T_93[34] ? 6'h22 : _ans_4_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_157 = _ans_4_leadingZeros_T_93[33] ? 6'h21 : _ans_4_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_158 = _ans_4_leadingZeros_T_93[32] ? 6'h20 : _ans_4_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_159 = _ans_4_leadingZeros_T_93[31] ? 6'h1f : _ans_4_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_160 = _ans_4_leadingZeros_T_93[30] ? 6'h1e : _ans_4_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_161 = _ans_4_leadingZeros_T_93[29] ? 6'h1d : _ans_4_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_162 = _ans_4_leadingZeros_T_93[28] ? 6'h1c : _ans_4_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_163 = _ans_4_leadingZeros_T_93[27] ? 6'h1b : _ans_4_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_164 = _ans_4_leadingZeros_T_93[26] ? 6'h1a : _ans_4_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_165 = _ans_4_leadingZeros_T_93[25] ? 6'h19 : _ans_4_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_166 = _ans_4_leadingZeros_T_93[24] ? 6'h18 : _ans_4_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_167 = _ans_4_leadingZeros_T_93[23] ? 6'h17 : _ans_4_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_168 = _ans_4_leadingZeros_T_93[22] ? 6'h16 : _ans_4_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_169 = _ans_4_leadingZeros_T_93[21] ? 6'h15 : _ans_4_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_170 = _ans_4_leadingZeros_T_93[20] ? 6'h14 : _ans_4_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_171 = _ans_4_leadingZeros_T_93[19] ? 6'h13 : _ans_4_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_172 = _ans_4_leadingZeros_T_93[18] ? 6'h12 : _ans_4_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_173 = _ans_4_leadingZeros_T_93[17] ? 6'h11 : _ans_4_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_174 = _ans_4_leadingZeros_T_93[16] ? 6'h10 : _ans_4_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_175 = _ans_4_leadingZeros_T_93[15] ? 6'hf : _ans_4_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_176 = _ans_4_leadingZeros_T_93[14] ? 6'he : _ans_4_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_177 = _ans_4_leadingZeros_T_93[13] ? 6'hd : _ans_4_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_178 = _ans_4_leadingZeros_T_93[12] ? 6'hc : _ans_4_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_179 = _ans_4_leadingZeros_T_93[11] ? 6'hb : _ans_4_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_180 = _ans_4_leadingZeros_T_93[10] ? 6'ha : _ans_4_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_181 = _ans_4_leadingZeros_T_93[9] ? 6'h9 : _ans_4_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_182 = _ans_4_leadingZeros_T_93[8] ? 6'h8 : _ans_4_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_183 = _ans_4_leadingZeros_T_93[7] ? 6'h7 : _ans_4_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_184 = _ans_4_leadingZeros_T_93[6] ? 6'h6 : _ans_4_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_185 = _ans_4_leadingZeros_T_93[5] ? 6'h5 : _ans_4_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_186 = _ans_4_leadingZeros_T_93[4] ? 6'h4 : _ans_4_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_187 = _ans_4_leadingZeros_T_93[3] ? 6'h3 : _ans_4_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_188 = _ans_4_leadingZeros_T_93[2] ? 6'h2 : _ans_4_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_leadingZeros_T_189 = _ans_4_leadingZeros_T_93[1] ? 6'h1 : _ans_4_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_4_leadingZeros = _ans_4_leadingZeros_T_93[0] ? 6'h0 : _ans_4_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_4_expRaw_T_1 = 6'h1f - ans_4_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_4_expRaw = ans_4_isZero ? 6'h0 : _ans_4_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_4_shiftAmt_T_2 = ans_4_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_4_shiftAmt = ans_4_expRaw > 6'h3 ? _ans_4_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_4_mantissaRaw_T = ans_4_absClipped >> ans_4_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_4_mantissaRaw = _ans_4_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_4_mantissa = ans_4_expRaw >= 6'h3 ? ans_4_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_4_expAdjusted = ans_4_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_4_exp_T_4 = ans_4_expAdjusted > 7'hf ? 4'hf : ans_4_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_4_exp = ans_4_isZero ? 4'h0 : _ans_4_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_4_fp8 = {ans_4_clippedX[31],ans_4_exp,ans_4_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_5 = {24'h0,linear_bias_5}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_5 = tempSum_5 + biasExtended_5; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_5_sign = sum32_5[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_5_absX_T = ~sum32_5; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_5_absX_T_2 = _ans_5_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_5_absX = ans_5_sign ? _ans_5_absX_T_2 : sum32_5; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_5_shiftedX_T_1 = _GEN_14432 - ans_5_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_5_shiftedX_T_3 = ans_5_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_5_shiftedX = ans_5_sign ? _ans_5_shiftedX_T_1 : _ans_5_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_5_scaledX_T_1 = ans_5_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_5_scaledX = _ans_5_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_5_clippedX_T_2 = ans_5_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_5_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_5_clippedX = ans_5_scaledX > 49'h1c0 ? 49'h1c0 : _ans_5_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_5_absClipped_T_1 = ~ans_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_5_absClipped_T_3 = _ans_5_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_5_absClipped = ans_5_clippedX[31] ? _ans_5_absClipped_T_3 : ans_5_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_5_isZero = ans_5_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39769 = {{16'd0}, ans_5_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_4 = _GEN_39769 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_6 = {ans_5_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_8 = _ans_5_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_9 = _ans_5_leadingZeros_T_4 | _ans_5_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39770 = {{8'd0}, _ans_5_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_14 = _GEN_39770 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_16 = {_ans_5_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_18 = _ans_5_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_19 = _ans_5_leadingZeros_T_14 | _ans_5_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39771 = {{4'd0}, _ans_5_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_24 = _GEN_39771 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_26 = {_ans_5_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_28 = _ans_5_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_29 = _ans_5_leadingZeros_T_24 | _ans_5_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39772 = {{2'd0}, _ans_5_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_34 = _GEN_39772 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_36 = {_ans_5_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_38 = _ans_5_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_39 = _ans_5_leadingZeros_T_34 | _ans_5_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39773 = {{1'd0}, _ans_5_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_44 = _GEN_39773 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_46 = {_ans_5_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_48 = _ans_5_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_5_leadingZeros_T_49 = _ans_5_leadingZeros_T_44 | _ans_5_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39774 = {{8'd0}, ans_5_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_55 = _GEN_39774 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_57 = {ans_5_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_59 = _ans_5_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_60 = _ans_5_leadingZeros_T_55 | _ans_5_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39775 = {{4'd0}, _ans_5_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_65 = _GEN_39775 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_67 = {_ans_5_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_69 = _ans_5_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_70 = _ans_5_leadingZeros_T_65 | _ans_5_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39776 = {{2'd0}, _ans_5_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_75 = _GEN_39776 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_77 = {_ans_5_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_79 = _ans_5_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_80 = _ans_5_leadingZeros_T_75 | _ans_5_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39777 = {{1'd0}, _ans_5_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_85 = _GEN_39777 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_87 = {_ans_5_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_89 = _ans_5_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_5_leadingZeros_T_90 = _ans_5_leadingZeros_T_85 | _ans_5_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_5_leadingZeros_T_93 = {_ans_5_leadingZeros_T_49,_ans_5_leadingZeros_T_90,ans_5_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_5_leadingZeros_T_143 = _ans_5_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_144 = _ans_5_leadingZeros_T_93[46] ? 6'h2e : _ans_5_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_145 = _ans_5_leadingZeros_T_93[45] ? 6'h2d : _ans_5_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_146 = _ans_5_leadingZeros_T_93[44] ? 6'h2c : _ans_5_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_147 = _ans_5_leadingZeros_T_93[43] ? 6'h2b : _ans_5_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_148 = _ans_5_leadingZeros_T_93[42] ? 6'h2a : _ans_5_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_149 = _ans_5_leadingZeros_T_93[41] ? 6'h29 : _ans_5_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_150 = _ans_5_leadingZeros_T_93[40] ? 6'h28 : _ans_5_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_151 = _ans_5_leadingZeros_T_93[39] ? 6'h27 : _ans_5_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_152 = _ans_5_leadingZeros_T_93[38] ? 6'h26 : _ans_5_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_153 = _ans_5_leadingZeros_T_93[37] ? 6'h25 : _ans_5_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_154 = _ans_5_leadingZeros_T_93[36] ? 6'h24 : _ans_5_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_155 = _ans_5_leadingZeros_T_93[35] ? 6'h23 : _ans_5_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_156 = _ans_5_leadingZeros_T_93[34] ? 6'h22 : _ans_5_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_157 = _ans_5_leadingZeros_T_93[33] ? 6'h21 : _ans_5_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_158 = _ans_5_leadingZeros_T_93[32] ? 6'h20 : _ans_5_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_159 = _ans_5_leadingZeros_T_93[31] ? 6'h1f : _ans_5_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_160 = _ans_5_leadingZeros_T_93[30] ? 6'h1e : _ans_5_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_161 = _ans_5_leadingZeros_T_93[29] ? 6'h1d : _ans_5_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_162 = _ans_5_leadingZeros_T_93[28] ? 6'h1c : _ans_5_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_163 = _ans_5_leadingZeros_T_93[27] ? 6'h1b : _ans_5_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_164 = _ans_5_leadingZeros_T_93[26] ? 6'h1a : _ans_5_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_165 = _ans_5_leadingZeros_T_93[25] ? 6'h19 : _ans_5_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_166 = _ans_5_leadingZeros_T_93[24] ? 6'h18 : _ans_5_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_167 = _ans_5_leadingZeros_T_93[23] ? 6'h17 : _ans_5_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_168 = _ans_5_leadingZeros_T_93[22] ? 6'h16 : _ans_5_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_169 = _ans_5_leadingZeros_T_93[21] ? 6'h15 : _ans_5_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_170 = _ans_5_leadingZeros_T_93[20] ? 6'h14 : _ans_5_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_171 = _ans_5_leadingZeros_T_93[19] ? 6'h13 : _ans_5_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_172 = _ans_5_leadingZeros_T_93[18] ? 6'h12 : _ans_5_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_173 = _ans_5_leadingZeros_T_93[17] ? 6'h11 : _ans_5_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_174 = _ans_5_leadingZeros_T_93[16] ? 6'h10 : _ans_5_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_175 = _ans_5_leadingZeros_T_93[15] ? 6'hf : _ans_5_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_176 = _ans_5_leadingZeros_T_93[14] ? 6'he : _ans_5_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_177 = _ans_5_leadingZeros_T_93[13] ? 6'hd : _ans_5_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_178 = _ans_5_leadingZeros_T_93[12] ? 6'hc : _ans_5_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_179 = _ans_5_leadingZeros_T_93[11] ? 6'hb : _ans_5_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_180 = _ans_5_leadingZeros_T_93[10] ? 6'ha : _ans_5_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_181 = _ans_5_leadingZeros_T_93[9] ? 6'h9 : _ans_5_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_182 = _ans_5_leadingZeros_T_93[8] ? 6'h8 : _ans_5_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_183 = _ans_5_leadingZeros_T_93[7] ? 6'h7 : _ans_5_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_184 = _ans_5_leadingZeros_T_93[6] ? 6'h6 : _ans_5_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_185 = _ans_5_leadingZeros_T_93[5] ? 6'h5 : _ans_5_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_186 = _ans_5_leadingZeros_T_93[4] ? 6'h4 : _ans_5_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_187 = _ans_5_leadingZeros_T_93[3] ? 6'h3 : _ans_5_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_188 = _ans_5_leadingZeros_T_93[2] ? 6'h2 : _ans_5_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_leadingZeros_T_189 = _ans_5_leadingZeros_T_93[1] ? 6'h1 : _ans_5_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_5_leadingZeros = _ans_5_leadingZeros_T_93[0] ? 6'h0 : _ans_5_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_5_expRaw_T_1 = 6'h1f - ans_5_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_5_expRaw = ans_5_isZero ? 6'h0 : _ans_5_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_5_shiftAmt_T_2 = ans_5_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_5_shiftAmt = ans_5_expRaw > 6'h3 ? _ans_5_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_5_mantissaRaw_T = ans_5_absClipped >> ans_5_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_5_mantissaRaw = _ans_5_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_5_mantissa = ans_5_expRaw >= 6'h3 ? ans_5_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_5_expAdjusted = ans_5_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_5_exp_T_4 = ans_5_expAdjusted > 7'hf ? 4'hf : ans_5_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_5_exp = ans_5_isZero ? 4'h0 : _ans_5_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_5_fp8 = {ans_5_clippedX[31],ans_5_exp,ans_5_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_6 = {24'h0,linear_bias_6}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_6 = tempSum_6 + biasExtended_6; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_6_sign = sum32_6[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_6_absX_T = ~sum32_6; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_6_absX_T_2 = _ans_6_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_6_absX = ans_6_sign ? _ans_6_absX_T_2 : sum32_6; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_6_shiftedX_T_1 = _GEN_14432 - ans_6_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_6_shiftedX_T_3 = ans_6_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_6_shiftedX = ans_6_sign ? _ans_6_shiftedX_T_1 : _ans_6_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_6_scaledX_T_1 = ans_6_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_6_scaledX = _ans_6_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_6_clippedX_T_2 = ans_6_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_6_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_6_clippedX = ans_6_scaledX > 49'h1c0 ? 49'h1c0 : _ans_6_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_6_absClipped_T_1 = ~ans_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_6_absClipped_T_3 = _ans_6_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_6_absClipped = ans_6_clippedX[31] ? _ans_6_absClipped_T_3 : ans_6_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_6_isZero = ans_6_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39780 = {{16'd0}, ans_6_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_4 = _GEN_39780 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_6 = {ans_6_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_8 = _ans_6_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_9 = _ans_6_leadingZeros_T_4 | _ans_6_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39781 = {{8'd0}, _ans_6_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_14 = _GEN_39781 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_16 = {_ans_6_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_18 = _ans_6_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_19 = _ans_6_leadingZeros_T_14 | _ans_6_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39782 = {{4'd0}, _ans_6_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_24 = _GEN_39782 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_26 = {_ans_6_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_28 = _ans_6_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_29 = _ans_6_leadingZeros_T_24 | _ans_6_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39783 = {{2'd0}, _ans_6_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_34 = _GEN_39783 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_36 = {_ans_6_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_38 = _ans_6_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_39 = _ans_6_leadingZeros_T_34 | _ans_6_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39784 = {{1'd0}, _ans_6_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_44 = _GEN_39784 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_46 = {_ans_6_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_48 = _ans_6_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_6_leadingZeros_T_49 = _ans_6_leadingZeros_T_44 | _ans_6_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39785 = {{8'd0}, ans_6_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_55 = _GEN_39785 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_57 = {ans_6_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_59 = _ans_6_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_60 = _ans_6_leadingZeros_T_55 | _ans_6_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39786 = {{4'd0}, _ans_6_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_65 = _GEN_39786 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_67 = {_ans_6_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_69 = _ans_6_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_70 = _ans_6_leadingZeros_T_65 | _ans_6_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39787 = {{2'd0}, _ans_6_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_75 = _GEN_39787 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_77 = {_ans_6_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_79 = _ans_6_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_80 = _ans_6_leadingZeros_T_75 | _ans_6_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39788 = {{1'd0}, _ans_6_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_85 = _GEN_39788 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_87 = {_ans_6_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_89 = _ans_6_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_6_leadingZeros_T_90 = _ans_6_leadingZeros_T_85 | _ans_6_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_6_leadingZeros_T_93 = {_ans_6_leadingZeros_T_49,_ans_6_leadingZeros_T_90,ans_6_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_6_leadingZeros_T_143 = _ans_6_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_144 = _ans_6_leadingZeros_T_93[46] ? 6'h2e : _ans_6_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_145 = _ans_6_leadingZeros_T_93[45] ? 6'h2d : _ans_6_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_146 = _ans_6_leadingZeros_T_93[44] ? 6'h2c : _ans_6_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_147 = _ans_6_leadingZeros_T_93[43] ? 6'h2b : _ans_6_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_148 = _ans_6_leadingZeros_T_93[42] ? 6'h2a : _ans_6_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_149 = _ans_6_leadingZeros_T_93[41] ? 6'h29 : _ans_6_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_150 = _ans_6_leadingZeros_T_93[40] ? 6'h28 : _ans_6_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_151 = _ans_6_leadingZeros_T_93[39] ? 6'h27 : _ans_6_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_152 = _ans_6_leadingZeros_T_93[38] ? 6'h26 : _ans_6_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_153 = _ans_6_leadingZeros_T_93[37] ? 6'h25 : _ans_6_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_154 = _ans_6_leadingZeros_T_93[36] ? 6'h24 : _ans_6_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_155 = _ans_6_leadingZeros_T_93[35] ? 6'h23 : _ans_6_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_156 = _ans_6_leadingZeros_T_93[34] ? 6'h22 : _ans_6_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_157 = _ans_6_leadingZeros_T_93[33] ? 6'h21 : _ans_6_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_158 = _ans_6_leadingZeros_T_93[32] ? 6'h20 : _ans_6_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_159 = _ans_6_leadingZeros_T_93[31] ? 6'h1f : _ans_6_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_160 = _ans_6_leadingZeros_T_93[30] ? 6'h1e : _ans_6_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_161 = _ans_6_leadingZeros_T_93[29] ? 6'h1d : _ans_6_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_162 = _ans_6_leadingZeros_T_93[28] ? 6'h1c : _ans_6_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_163 = _ans_6_leadingZeros_T_93[27] ? 6'h1b : _ans_6_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_164 = _ans_6_leadingZeros_T_93[26] ? 6'h1a : _ans_6_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_165 = _ans_6_leadingZeros_T_93[25] ? 6'h19 : _ans_6_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_166 = _ans_6_leadingZeros_T_93[24] ? 6'h18 : _ans_6_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_167 = _ans_6_leadingZeros_T_93[23] ? 6'h17 : _ans_6_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_168 = _ans_6_leadingZeros_T_93[22] ? 6'h16 : _ans_6_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_169 = _ans_6_leadingZeros_T_93[21] ? 6'h15 : _ans_6_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_170 = _ans_6_leadingZeros_T_93[20] ? 6'h14 : _ans_6_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_171 = _ans_6_leadingZeros_T_93[19] ? 6'h13 : _ans_6_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_172 = _ans_6_leadingZeros_T_93[18] ? 6'h12 : _ans_6_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_173 = _ans_6_leadingZeros_T_93[17] ? 6'h11 : _ans_6_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_174 = _ans_6_leadingZeros_T_93[16] ? 6'h10 : _ans_6_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_175 = _ans_6_leadingZeros_T_93[15] ? 6'hf : _ans_6_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_176 = _ans_6_leadingZeros_T_93[14] ? 6'he : _ans_6_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_177 = _ans_6_leadingZeros_T_93[13] ? 6'hd : _ans_6_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_178 = _ans_6_leadingZeros_T_93[12] ? 6'hc : _ans_6_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_179 = _ans_6_leadingZeros_T_93[11] ? 6'hb : _ans_6_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_180 = _ans_6_leadingZeros_T_93[10] ? 6'ha : _ans_6_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_181 = _ans_6_leadingZeros_T_93[9] ? 6'h9 : _ans_6_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_182 = _ans_6_leadingZeros_T_93[8] ? 6'h8 : _ans_6_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_183 = _ans_6_leadingZeros_T_93[7] ? 6'h7 : _ans_6_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_184 = _ans_6_leadingZeros_T_93[6] ? 6'h6 : _ans_6_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_185 = _ans_6_leadingZeros_T_93[5] ? 6'h5 : _ans_6_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_186 = _ans_6_leadingZeros_T_93[4] ? 6'h4 : _ans_6_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_187 = _ans_6_leadingZeros_T_93[3] ? 6'h3 : _ans_6_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_188 = _ans_6_leadingZeros_T_93[2] ? 6'h2 : _ans_6_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_leadingZeros_T_189 = _ans_6_leadingZeros_T_93[1] ? 6'h1 : _ans_6_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_6_leadingZeros = _ans_6_leadingZeros_T_93[0] ? 6'h0 : _ans_6_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_6_expRaw_T_1 = 6'h1f - ans_6_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_6_expRaw = ans_6_isZero ? 6'h0 : _ans_6_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_6_shiftAmt_T_2 = ans_6_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_6_shiftAmt = ans_6_expRaw > 6'h3 ? _ans_6_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_6_mantissaRaw_T = ans_6_absClipped >> ans_6_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_6_mantissaRaw = _ans_6_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_6_mantissa = ans_6_expRaw >= 6'h3 ? ans_6_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_6_expAdjusted = ans_6_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_6_exp_T_4 = ans_6_expAdjusted > 7'hf ? 4'hf : ans_6_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_6_exp = ans_6_isZero ? 4'h0 : _ans_6_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_6_fp8 = {ans_6_clippedX[31],ans_6_exp,ans_6_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_7 = {24'h0,linear_bias_7}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_7 = tempSum_7 + biasExtended_7; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_7_sign = sum32_7[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_7_absX_T = ~sum32_7; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_7_absX_T_2 = _ans_7_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_7_absX = ans_7_sign ? _ans_7_absX_T_2 : sum32_7; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_7_shiftedX_T_1 = _GEN_14432 - ans_7_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_7_shiftedX_T_3 = ans_7_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_7_shiftedX = ans_7_sign ? _ans_7_shiftedX_T_1 : _ans_7_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_7_scaledX_T_1 = ans_7_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_7_scaledX = _ans_7_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_7_clippedX_T_2 = ans_7_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_7_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_7_clippedX = ans_7_scaledX > 49'h1c0 ? 49'h1c0 : _ans_7_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_7_absClipped_T_1 = ~ans_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_7_absClipped_T_3 = _ans_7_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_7_absClipped = ans_7_clippedX[31] ? _ans_7_absClipped_T_3 : ans_7_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_7_isZero = ans_7_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39791 = {{16'd0}, ans_7_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_4 = _GEN_39791 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_6 = {ans_7_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_8 = _ans_7_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_9 = _ans_7_leadingZeros_T_4 | _ans_7_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39792 = {{8'd0}, _ans_7_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_14 = _GEN_39792 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_16 = {_ans_7_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_18 = _ans_7_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_19 = _ans_7_leadingZeros_T_14 | _ans_7_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39793 = {{4'd0}, _ans_7_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_24 = _GEN_39793 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_26 = {_ans_7_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_28 = _ans_7_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_29 = _ans_7_leadingZeros_T_24 | _ans_7_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39794 = {{2'd0}, _ans_7_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_34 = _GEN_39794 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_36 = {_ans_7_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_38 = _ans_7_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_39 = _ans_7_leadingZeros_T_34 | _ans_7_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39795 = {{1'd0}, _ans_7_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_44 = _GEN_39795 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_46 = {_ans_7_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_48 = _ans_7_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_7_leadingZeros_T_49 = _ans_7_leadingZeros_T_44 | _ans_7_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39796 = {{8'd0}, ans_7_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_55 = _GEN_39796 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_57 = {ans_7_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_59 = _ans_7_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_60 = _ans_7_leadingZeros_T_55 | _ans_7_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39797 = {{4'd0}, _ans_7_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_65 = _GEN_39797 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_67 = {_ans_7_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_69 = _ans_7_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_70 = _ans_7_leadingZeros_T_65 | _ans_7_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39798 = {{2'd0}, _ans_7_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_75 = _GEN_39798 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_77 = {_ans_7_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_79 = _ans_7_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_80 = _ans_7_leadingZeros_T_75 | _ans_7_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39799 = {{1'd0}, _ans_7_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_85 = _GEN_39799 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_87 = {_ans_7_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_89 = _ans_7_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_7_leadingZeros_T_90 = _ans_7_leadingZeros_T_85 | _ans_7_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_7_leadingZeros_T_93 = {_ans_7_leadingZeros_T_49,_ans_7_leadingZeros_T_90,ans_7_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_7_leadingZeros_T_143 = _ans_7_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_144 = _ans_7_leadingZeros_T_93[46] ? 6'h2e : _ans_7_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_145 = _ans_7_leadingZeros_T_93[45] ? 6'h2d : _ans_7_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_146 = _ans_7_leadingZeros_T_93[44] ? 6'h2c : _ans_7_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_147 = _ans_7_leadingZeros_T_93[43] ? 6'h2b : _ans_7_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_148 = _ans_7_leadingZeros_T_93[42] ? 6'h2a : _ans_7_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_149 = _ans_7_leadingZeros_T_93[41] ? 6'h29 : _ans_7_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_150 = _ans_7_leadingZeros_T_93[40] ? 6'h28 : _ans_7_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_151 = _ans_7_leadingZeros_T_93[39] ? 6'h27 : _ans_7_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_152 = _ans_7_leadingZeros_T_93[38] ? 6'h26 : _ans_7_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_153 = _ans_7_leadingZeros_T_93[37] ? 6'h25 : _ans_7_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_154 = _ans_7_leadingZeros_T_93[36] ? 6'h24 : _ans_7_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_155 = _ans_7_leadingZeros_T_93[35] ? 6'h23 : _ans_7_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_156 = _ans_7_leadingZeros_T_93[34] ? 6'h22 : _ans_7_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_157 = _ans_7_leadingZeros_T_93[33] ? 6'h21 : _ans_7_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_158 = _ans_7_leadingZeros_T_93[32] ? 6'h20 : _ans_7_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_159 = _ans_7_leadingZeros_T_93[31] ? 6'h1f : _ans_7_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_160 = _ans_7_leadingZeros_T_93[30] ? 6'h1e : _ans_7_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_161 = _ans_7_leadingZeros_T_93[29] ? 6'h1d : _ans_7_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_162 = _ans_7_leadingZeros_T_93[28] ? 6'h1c : _ans_7_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_163 = _ans_7_leadingZeros_T_93[27] ? 6'h1b : _ans_7_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_164 = _ans_7_leadingZeros_T_93[26] ? 6'h1a : _ans_7_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_165 = _ans_7_leadingZeros_T_93[25] ? 6'h19 : _ans_7_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_166 = _ans_7_leadingZeros_T_93[24] ? 6'h18 : _ans_7_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_167 = _ans_7_leadingZeros_T_93[23] ? 6'h17 : _ans_7_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_168 = _ans_7_leadingZeros_T_93[22] ? 6'h16 : _ans_7_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_169 = _ans_7_leadingZeros_T_93[21] ? 6'h15 : _ans_7_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_170 = _ans_7_leadingZeros_T_93[20] ? 6'h14 : _ans_7_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_171 = _ans_7_leadingZeros_T_93[19] ? 6'h13 : _ans_7_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_172 = _ans_7_leadingZeros_T_93[18] ? 6'h12 : _ans_7_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_173 = _ans_7_leadingZeros_T_93[17] ? 6'h11 : _ans_7_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_174 = _ans_7_leadingZeros_T_93[16] ? 6'h10 : _ans_7_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_175 = _ans_7_leadingZeros_T_93[15] ? 6'hf : _ans_7_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_176 = _ans_7_leadingZeros_T_93[14] ? 6'he : _ans_7_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_177 = _ans_7_leadingZeros_T_93[13] ? 6'hd : _ans_7_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_178 = _ans_7_leadingZeros_T_93[12] ? 6'hc : _ans_7_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_179 = _ans_7_leadingZeros_T_93[11] ? 6'hb : _ans_7_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_180 = _ans_7_leadingZeros_T_93[10] ? 6'ha : _ans_7_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_181 = _ans_7_leadingZeros_T_93[9] ? 6'h9 : _ans_7_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_182 = _ans_7_leadingZeros_T_93[8] ? 6'h8 : _ans_7_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_183 = _ans_7_leadingZeros_T_93[7] ? 6'h7 : _ans_7_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_184 = _ans_7_leadingZeros_T_93[6] ? 6'h6 : _ans_7_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_185 = _ans_7_leadingZeros_T_93[5] ? 6'h5 : _ans_7_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_186 = _ans_7_leadingZeros_T_93[4] ? 6'h4 : _ans_7_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_187 = _ans_7_leadingZeros_T_93[3] ? 6'h3 : _ans_7_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_188 = _ans_7_leadingZeros_T_93[2] ? 6'h2 : _ans_7_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_leadingZeros_T_189 = _ans_7_leadingZeros_T_93[1] ? 6'h1 : _ans_7_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_7_leadingZeros = _ans_7_leadingZeros_T_93[0] ? 6'h0 : _ans_7_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_7_expRaw_T_1 = 6'h1f - ans_7_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_7_expRaw = ans_7_isZero ? 6'h0 : _ans_7_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_7_shiftAmt_T_2 = ans_7_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_7_shiftAmt = ans_7_expRaw > 6'h3 ? _ans_7_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_7_mantissaRaw_T = ans_7_absClipped >> ans_7_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_7_mantissaRaw = _ans_7_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_7_mantissa = ans_7_expRaw >= 6'h3 ? ans_7_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_7_expAdjusted = ans_7_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_7_exp_T_4 = ans_7_expAdjusted > 7'hf ? 4'hf : ans_7_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_7_exp = ans_7_isZero ? 4'h0 : _ans_7_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_7_fp8 = {ans_7_clippedX[31],ans_7_exp,ans_7_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_8 = {24'h0,linear_bias_8}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_8 = tempSum_8 + biasExtended_8; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_8_sign = sum32_8[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_8_absX_T = ~sum32_8; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_8_absX_T_2 = _ans_8_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_8_absX = ans_8_sign ? _ans_8_absX_T_2 : sum32_8; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_8_shiftedX_T_1 = _GEN_14432 - ans_8_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_8_shiftedX_T_3 = ans_8_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_8_shiftedX = ans_8_sign ? _ans_8_shiftedX_T_1 : _ans_8_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_8_scaledX_T_1 = ans_8_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_8_scaledX = _ans_8_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_8_clippedX_T_2 = ans_8_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_8_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_8_clippedX = ans_8_scaledX > 49'h1c0 ? 49'h1c0 : _ans_8_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_8_absClipped_T_1 = ~ans_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_8_absClipped_T_3 = _ans_8_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_8_absClipped = ans_8_clippedX[31] ? _ans_8_absClipped_T_3 : ans_8_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_8_isZero = ans_8_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39802 = {{16'd0}, ans_8_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_4 = _GEN_39802 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_6 = {ans_8_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_8 = _ans_8_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_9 = _ans_8_leadingZeros_T_4 | _ans_8_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39803 = {{8'd0}, _ans_8_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_14 = _GEN_39803 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_16 = {_ans_8_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_18 = _ans_8_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_19 = _ans_8_leadingZeros_T_14 | _ans_8_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39804 = {{4'd0}, _ans_8_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_24 = _GEN_39804 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_26 = {_ans_8_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_28 = _ans_8_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_29 = _ans_8_leadingZeros_T_24 | _ans_8_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39805 = {{2'd0}, _ans_8_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_34 = _GEN_39805 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_36 = {_ans_8_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_38 = _ans_8_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_39 = _ans_8_leadingZeros_T_34 | _ans_8_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39806 = {{1'd0}, _ans_8_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_44 = _GEN_39806 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_46 = {_ans_8_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_48 = _ans_8_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_8_leadingZeros_T_49 = _ans_8_leadingZeros_T_44 | _ans_8_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39807 = {{8'd0}, ans_8_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_55 = _GEN_39807 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_57 = {ans_8_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_59 = _ans_8_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_60 = _ans_8_leadingZeros_T_55 | _ans_8_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39808 = {{4'd0}, _ans_8_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_65 = _GEN_39808 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_67 = {_ans_8_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_69 = _ans_8_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_70 = _ans_8_leadingZeros_T_65 | _ans_8_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39809 = {{2'd0}, _ans_8_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_75 = _GEN_39809 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_77 = {_ans_8_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_79 = _ans_8_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_80 = _ans_8_leadingZeros_T_75 | _ans_8_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39810 = {{1'd0}, _ans_8_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_85 = _GEN_39810 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_87 = {_ans_8_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_89 = _ans_8_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_8_leadingZeros_T_90 = _ans_8_leadingZeros_T_85 | _ans_8_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_8_leadingZeros_T_93 = {_ans_8_leadingZeros_T_49,_ans_8_leadingZeros_T_90,ans_8_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_8_leadingZeros_T_143 = _ans_8_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_144 = _ans_8_leadingZeros_T_93[46] ? 6'h2e : _ans_8_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_145 = _ans_8_leadingZeros_T_93[45] ? 6'h2d : _ans_8_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_146 = _ans_8_leadingZeros_T_93[44] ? 6'h2c : _ans_8_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_147 = _ans_8_leadingZeros_T_93[43] ? 6'h2b : _ans_8_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_148 = _ans_8_leadingZeros_T_93[42] ? 6'h2a : _ans_8_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_149 = _ans_8_leadingZeros_T_93[41] ? 6'h29 : _ans_8_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_150 = _ans_8_leadingZeros_T_93[40] ? 6'h28 : _ans_8_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_151 = _ans_8_leadingZeros_T_93[39] ? 6'h27 : _ans_8_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_152 = _ans_8_leadingZeros_T_93[38] ? 6'h26 : _ans_8_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_153 = _ans_8_leadingZeros_T_93[37] ? 6'h25 : _ans_8_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_154 = _ans_8_leadingZeros_T_93[36] ? 6'h24 : _ans_8_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_155 = _ans_8_leadingZeros_T_93[35] ? 6'h23 : _ans_8_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_156 = _ans_8_leadingZeros_T_93[34] ? 6'h22 : _ans_8_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_157 = _ans_8_leadingZeros_T_93[33] ? 6'h21 : _ans_8_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_158 = _ans_8_leadingZeros_T_93[32] ? 6'h20 : _ans_8_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_159 = _ans_8_leadingZeros_T_93[31] ? 6'h1f : _ans_8_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_160 = _ans_8_leadingZeros_T_93[30] ? 6'h1e : _ans_8_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_161 = _ans_8_leadingZeros_T_93[29] ? 6'h1d : _ans_8_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_162 = _ans_8_leadingZeros_T_93[28] ? 6'h1c : _ans_8_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_163 = _ans_8_leadingZeros_T_93[27] ? 6'h1b : _ans_8_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_164 = _ans_8_leadingZeros_T_93[26] ? 6'h1a : _ans_8_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_165 = _ans_8_leadingZeros_T_93[25] ? 6'h19 : _ans_8_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_166 = _ans_8_leadingZeros_T_93[24] ? 6'h18 : _ans_8_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_167 = _ans_8_leadingZeros_T_93[23] ? 6'h17 : _ans_8_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_168 = _ans_8_leadingZeros_T_93[22] ? 6'h16 : _ans_8_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_169 = _ans_8_leadingZeros_T_93[21] ? 6'h15 : _ans_8_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_170 = _ans_8_leadingZeros_T_93[20] ? 6'h14 : _ans_8_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_171 = _ans_8_leadingZeros_T_93[19] ? 6'h13 : _ans_8_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_172 = _ans_8_leadingZeros_T_93[18] ? 6'h12 : _ans_8_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_173 = _ans_8_leadingZeros_T_93[17] ? 6'h11 : _ans_8_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_174 = _ans_8_leadingZeros_T_93[16] ? 6'h10 : _ans_8_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_175 = _ans_8_leadingZeros_T_93[15] ? 6'hf : _ans_8_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_176 = _ans_8_leadingZeros_T_93[14] ? 6'he : _ans_8_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_177 = _ans_8_leadingZeros_T_93[13] ? 6'hd : _ans_8_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_178 = _ans_8_leadingZeros_T_93[12] ? 6'hc : _ans_8_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_179 = _ans_8_leadingZeros_T_93[11] ? 6'hb : _ans_8_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_180 = _ans_8_leadingZeros_T_93[10] ? 6'ha : _ans_8_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_181 = _ans_8_leadingZeros_T_93[9] ? 6'h9 : _ans_8_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_182 = _ans_8_leadingZeros_T_93[8] ? 6'h8 : _ans_8_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_183 = _ans_8_leadingZeros_T_93[7] ? 6'h7 : _ans_8_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_184 = _ans_8_leadingZeros_T_93[6] ? 6'h6 : _ans_8_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_185 = _ans_8_leadingZeros_T_93[5] ? 6'h5 : _ans_8_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_186 = _ans_8_leadingZeros_T_93[4] ? 6'h4 : _ans_8_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_187 = _ans_8_leadingZeros_T_93[3] ? 6'h3 : _ans_8_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_188 = _ans_8_leadingZeros_T_93[2] ? 6'h2 : _ans_8_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_leadingZeros_T_189 = _ans_8_leadingZeros_T_93[1] ? 6'h1 : _ans_8_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_8_leadingZeros = _ans_8_leadingZeros_T_93[0] ? 6'h0 : _ans_8_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_8_expRaw_T_1 = 6'h1f - ans_8_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_8_expRaw = ans_8_isZero ? 6'h0 : _ans_8_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_8_shiftAmt_T_2 = ans_8_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_8_shiftAmt = ans_8_expRaw > 6'h3 ? _ans_8_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_8_mantissaRaw_T = ans_8_absClipped >> ans_8_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_8_mantissaRaw = _ans_8_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_8_mantissa = ans_8_expRaw >= 6'h3 ? ans_8_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_8_expAdjusted = ans_8_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_8_exp_T_4 = ans_8_expAdjusted > 7'hf ? 4'hf : ans_8_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_8_exp = ans_8_isZero ? 4'h0 : _ans_8_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_8_fp8 = {ans_8_clippedX[31],ans_8_exp,ans_8_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_9 = {24'h0,linear_bias_9}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_9 = tempSum_9 + biasExtended_9; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_9_sign = sum32_9[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_9_absX_T = ~sum32_9; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_9_absX_T_2 = _ans_9_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_9_absX = ans_9_sign ? _ans_9_absX_T_2 : sum32_9; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_9_shiftedX_T_1 = _GEN_14432 - ans_9_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_9_shiftedX_T_3 = ans_9_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_9_shiftedX = ans_9_sign ? _ans_9_shiftedX_T_1 : _ans_9_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_9_scaledX_T_1 = ans_9_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_9_scaledX = _ans_9_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_9_clippedX_T_2 = ans_9_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_9_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_9_clippedX = ans_9_scaledX > 49'h1c0 ? 49'h1c0 : _ans_9_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_9_absClipped_T_1 = ~ans_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_9_absClipped_T_3 = _ans_9_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_9_absClipped = ans_9_clippedX[31] ? _ans_9_absClipped_T_3 : ans_9_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_9_isZero = ans_9_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39813 = {{16'd0}, ans_9_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_4 = _GEN_39813 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_6 = {ans_9_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_8 = _ans_9_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_9 = _ans_9_leadingZeros_T_4 | _ans_9_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39814 = {{8'd0}, _ans_9_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_14 = _GEN_39814 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_16 = {_ans_9_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_18 = _ans_9_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_19 = _ans_9_leadingZeros_T_14 | _ans_9_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39815 = {{4'd0}, _ans_9_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_24 = _GEN_39815 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_26 = {_ans_9_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_28 = _ans_9_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_29 = _ans_9_leadingZeros_T_24 | _ans_9_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39816 = {{2'd0}, _ans_9_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_34 = _GEN_39816 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_36 = {_ans_9_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_38 = _ans_9_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_39 = _ans_9_leadingZeros_T_34 | _ans_9_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39817 = {{1'd0}, _ans_9_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_44 = _GEN_39817 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_46 = {_ans_9_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_48 = _ans_9_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_9_leadingZeros_T_49 = _ans_9_leadingZeros_T_44 | _ans_9_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39818 = {{8'd0}, ans_9_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_55 = _GEN_39818 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_57 = {ans_9_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_59 = _ans_9_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_60 = _ans_9_leadingZeros_T_55 | _ans_9_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39819 = {{4'd0}, _ans_9_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_65 = _GEN_39819 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_67 = {_ans_9_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_69 = _ans_9_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_70 = _ans_9_leadingZeros_T_65 | _ans_9_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39820 = {{2'd0}, _ans_9_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_75 = _GEN_39820 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_77 = {_ans_9_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_79 = _ans_9_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_80 = _ans_9_leadingZeros_T_75 | _ans_9_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39821 = {{1'd0}, _ans_9_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_85 = _GEN_39821 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_87 = {_ans_9_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_89 = _ans_9_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_9_leadingZeros_T_90 = _ans_9_leadingZeros_T_85 | _ans_9_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_9_leadingZeros_T_93 = {_ans_9_leadingZeros_T_49,_ans_9_leadingZeros_T_90,ans_9_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_9_leadingZeros_T_143 = _ans_9_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_144 = _ans_9_leadingZeros_T_93[46] ? 6'h2e : _ans_9_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_145 = _ans_9_leadingZeros_T_93[45] ? 6'h2d : _ans_9_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_146 = _ans_9_leadingZeros_T_93[44] ? 6'h2c : _ans_9_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_147 = _ans_9_leadingZeros_T_93[43] ? 6'h2b : _ans_9_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_148 = _ans_9_leadingZeros_T_93[42] ? 6'h2a : _ans_9_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_149 = _ans_9_leadingZeros_T_93[41] ? 6'h29 : _ans_9_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_150 = _ans_9_leadingZeros_T_93[40] ? 6'h28 : _ans_9_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_151 = _ans_9_leadingZeros_T_93[39] ? 6'h27 : _ans_9_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_152 = _ans_9_leadingZeros_T_93[38] ? 6'h26 : _ans_9_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_153 = _ans_9_leadingZeros_T_93[37] ? 6'h25 : _ans_9_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_154 = _ans_9_leadingZeros_T_93[36] ? 6'h24 : _ans_9_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_155 = _ans_9_leadingZeros_T_93[35] ? 6'h23 : _ans_9_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_156 = _ans_9_leadingZeros_T_93[34] ? 6'h22 : _ans_9_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_157 = _ans_9_leadingZeros_T_93[33] ? 6'h21 : _ans_9_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_158 = _ans_9_leadingZeros_T_93[32] ? 6'h20 : _ans_9_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_159 = _ans_9_leadingZeros_T_93[31] ? 6'h1f : _ans_9_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_160 = _ans_9_leadingZeros_T_93[30] ? 6'h1e : _ans_9_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_161 = _ans_9_leadingZeros_T_93[29] ? 6'h1d : _ans_9_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_162 = _ans_9_leadingZeros_T_93[28] ? 6'h1c : _ans_9_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_163 = _ans_9_leadingZeros_T_93[27] ? 6'h1b : _ans_9_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_164 = _ans_9_leadingZeros_T_93[26] ? 6'h1a : _ans_9_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_165 = _ans_9_leadingZeros_T_93[25] ? 6'h19 : _ans_9_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_166 = _ans_9_leadingZeros_T_93[24] ? 6'h18 : _ans_9_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_167 = _ans_9_leadingZeros_T_93[23] ? 6'h17 : _ans_9_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_168 = _ans_9_leadingZeros_T_93[22] ? 6'h16 : _ans_9_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_169 = _ans_9_leadingZeros_T_93[21] ? 6'h15 : _ans_9_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_170 = _ans_9_leadingZeros_T_93[20] ? 6'h14 : _ans_9_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_171 = _ans_9_leadingZeros_T_93[19] ? 6'h13 : _ans_9_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_172 = _ans_9_leadingZeros_T_93[18] ? 6'h12 : _ans_9_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_173 = _ans_9_leadingZeros_T_93[17] ? 6'h11 : _ans_9_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_174 = _ans_9_leadingZeros_T_93[16] ? 6'h10 : _ans_9_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_175 = _ans_9_leadingZeros_T_93[15] ? 6'hf : _ans_9_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_176 = _ans_9_leadingZeros_T_93[14] ? 6'he : _ans_9_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_177 = _ans_9_leadingZeros_T_93[13] ? 6'hd : _ans_9_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_178 = _ans_9_leadingZeros_T_93[12] ? 6'hc : _ans_9_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_179 = _ans_9_leadingZeros_T_93[11] ? 6'hb : _ans_9_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_180 = _ans_9_leadingZeros_T_93[10] ? 6'ha : _ans_9_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_181 = _ans_9_leadingZeros_T_93[9] ? 6'h9 : _ans_9_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_182 = _ans_9_leadingZeros_T_93[8] ? 6'h8 : _ans_9_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_183 = _ans_9_leadingZeros_T_93[7] ? 6'h7 : _ans_9_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_184 = _ans_9_leadingZeros_T_93[6] ? 6'h6 : _ans_9_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_185 = _ans_9_leadingZeros_T_93[5] ? 6'h5 : _ans_9_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_186 = _ans_9_leadingZeros_T_93[4] ? 6'h4 : _ans_9_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_187 = _ans_9_leadingZeros_T_93[3] ? 6'h3 : _ans_9_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_188 = _ans_9_leadingZeros_T_93[2] ? 6'h2 : _ans_9_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_leadingZeros_T_189 = _ans_9_leadingZeros_T_93[1] ? 6'h1 : _ans_9_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_9_leadingZeros = _ans_9_leadingZeros_T_93[0] ? 6'h0 : _ans_9_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_9_expRaw_T_1 = 6'h1f - ans_9_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_9_expRaw = ans_9_isZero ? 6'h0 : _ans_9_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_9_shiftAmt_T_2 = ans_9_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_9_shiftAmt = ans_9_expRaw > 6'h3 ? _ans_9_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_9_mantissaRaw_T = ans_9_absClipped >> ans_9_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_9_mantissaRaw = _ans_9_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_9_mantissa = ans_9_expRaw >= 6'h3 ? ans_9_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_9_expAdjusted = ans_9_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_9_exp_T_4 = ans_9_expAdjusted > 7'hf ? 4'hf : ans_9_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_9_exp = ans_9_isZero ? 4'h0 : _ans_9_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_9_fp8 = {ans_9_clippedX[31],ans_9_exp,ans_9_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_10 = {24'h0,linear_bias_10}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_10 = tempSum_10 + biasExtended_10; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_10_sign = sum32_10[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_10_absX_T = ~sum32_10; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_10_absX_T_2 = _ans_10_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_10_absX = ans_10_sign ? _ans_10_absX_T_2 : sum32_10; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_10_shiftedX_T_1 = _GEN_14432 - ans_10_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_10_shiftedX_T_3 = ans_10_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_10_shiftedX = ans_10_sign ? _ans_10_shiftedX_T_1 : _ans_10_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_10_scaledX_T_1 = ans_10_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_10_scaledX = _ans_10_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_10_clippedX_T_2 = ans_10_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_10_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_10_clippedX = ans_10_scaledX > 49'h1c0 ? 49'h1c0 : _ans_10_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_10_absClipped_T_1 = ~ans_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_10_absClipped_T_3 = _ans_10_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_10_absClipped = ans_10_clippedX[31] ? _ans_10_absClipped_T_3 : ans_10_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_10_isZero = ans_10_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39824 = {{16'd0}, ans_10_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_4 = _GEN_39824 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_6 = {ans_10_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_8 = _ans_10_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_9 = _ans_10_leadingZeros_T_4 | _ans_10_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39825 = {{8'd0}, _ans_10_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_14 = _GEN_39825 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_16 = {_ans_10_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_18 = _ans_10_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_19 = _ans_10_leadingZeros_T_14 | _ans_10_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39826 = {{4'd0}, _ans_10_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_24 = _GEN_39826 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_26 = {_ans_10_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_28 = _ans_10_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_29 = _ans_10_leadingZeros_T_24 | _ans_10_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39827 = {{2'd0}, _ans_10_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_34 = _GEN_39827 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_36 = {_ans_10_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_38 = _ans_10_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_39 = _ans_10_leadingZeros_T_34 | _ans_10_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39828 = {{1'd0}, _ans_10_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_44 = _GEN_39828 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_46 = {_ans_10_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_48 = _ans_10_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_10_leadingZeros_T_49 = _ans_10_leadingZeros_T_44 | _ans_10_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39829 = {{8'd0}, ans_10_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_55 = _GEN_39829 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_57 = {ans_10_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_59 = _ans_10_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_60 = _ans_10_leadingZeros_T_55 | _ans_10_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39830 = {{4'd0}, _ans_10_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_65 = _GEN_39830 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_67 = {_ans_10_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_69 = _ans_10_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_70 = _ans_10_leadingZeros_T_65 | _ans_10_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39831 = {{2'd0}, _ans_10_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_75 = _GEN_39831 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_77 = {_ans_10_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_79 = _ans_10_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_80 = _ans_10_leadingZeros_T_75 | _ans_10_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39832 = {{1'd0}, _ans_10_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_85 = _GEN_39832 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_87 = {_ans_10_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_89 = _ans_10_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_10_leadingZeros_T_90 = _ans_10_leadingZeros_T_85 | _ans_10_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_10_leadingZeros_T_93 = {_ans_10_leadingZeros_T_49,_ans_10_leadingZeros_T_90,ans_10_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_10_leadingZeros_T_143 = _ans_10_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_144 = _ans_10_leadingZeros_T_93[46] ? 6'h2e : _ans_10_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_145 = _ans_10_leadingZeros_T_93[45] ? 6'h2d : _ans_10_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_146 = _ans_10_leadingZeros_T_93[44] ? 6'h2c : _ans_10_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_147 = _ans_10_leadingZeros_T_93[43] ? 6'h2b : _ans_10_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_148 = _ans_10_leadingZeros_T_93[42] ? 6'h2a : _ans_10_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_149 = _ans_10_leadingZeros_T_93[41] ? 6'h29 : _ans_10_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_150 = _ans_10_leadingZeros_T_93[40] ? 6'h28 : _ans_10_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_151 = _ans_10_leadingZeros_T_93[39] ? 6'h27 : _ans_10_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_152 = _ans_10_leadingZeros_T_93[38] ? 6'h26 : _ans_10_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_153 = _ans_10_leadingZeros_T_93[37] ? 6'h25 : _ans_10_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_154 = _ans_10_leadingZeros_T_93[36] ? 6'h24 : _ans_10_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_155 = _ans_10_leadingZeros_T_93[35] ? 6'h23 : _ans_10_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_156 = _ans_10_leadingZeros_T_93[34] ? 6'h22 : _ans_10_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_157 = _ans_10_leadingZeros_T_93[33] ? 6'h21 : _ans_10_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_158 = _ans_10_leadingZeros_T_93[32] ? 6'h20 : _ans_10_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_159 = _ans_10_leadingZeros_T_93[31] ? 6'h1f : _ans_10_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_160 = _ans_10_leadingZeros_T_93[30] ? 6'h1e : _ans_10_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_161 = _ans_10_leadingZeros_T_93[29] ? 6'h1d : _ans_10_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_162 = _ans_10_leadingZeros_T_93[28] ? 6'h1c : _ans_10_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_163 = _ans_10_leadingZeros_T_93[27] ? 6'h1b : _ans_10_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_164 = _ans_10_leadingZeros_T_93[26] ? 6'h1a : _ans_10_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_165 = _ans_10_leadingZeros_T_93[25] ? 6'h19 : _ans_10_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_166 = _ans_10_leadingZeros_T_93[24] ? 6'h18 : _ans_10_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_167 = _ans_10_leadingZeros_T_93[23] ? 6'h17 : _ans_10_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_168 = _ans_10_leadingZeros_T_93[22] ? 6'h16 : _ans_10_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_169 = _ans_10_leadingZeros_T_93[21] ? 6'h15 : _ans_10_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_170 = _ans_10_leadingZeros_T_93[20] ? 6'h14 : _ans_10_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_171 = _ans_10_leadingZeros_T_93[19] ? 6'h13 : _ans_10_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_172 = _ans_10_leadingZeros_T_93[18] ? 6'h12 : _ans_10_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_173 = _ans_10_leadingZeros_T_93[17] ? 6'h11 : _ans_10_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_174 = _ans_10_leadingZeros_T_93[16] ? 6'h10 : _ans_10_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_175 = _ans_10_leadingZeros_T_93[15] ? 6'hf : _ans_10_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_176 = _ans_10_leadingZeros_T_93[14] ? 6'he : _ans_10_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_177 = _ans_10_leadingZeros_T_93[13] ? 6'hd : _ans_10_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_178 = _ans_10_leadingZeros_T_93[12] ? 6'hc : _ans_10_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_179 = _ans_10_leadingZeros_T_93[11] ? 6'hb : _ans_10_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_180 = _ans_10_leadingZeros_T_93[10] ? 6'ha : _ans_10_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_181 = _ans_10_leadingZeros_T_93[9] ? 6'h9 : _ans_10_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_182 = _ans_10_leadingZeros_T_93[8] ? 6'h8 : _ans_10_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_183 = _ans_10_leadingZeros_T_93[7] ? 6'h7 : _ans_10_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_184 = _ans_10_leadingZeros_T_93[6] ? 6'h6 : _ans_10_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_185 = _ans_10_leadingZeros_T_93[5] ? 6'h5 : _ans_10_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_186 = _ans_10_leadingZeros_T_93[4] ? 6'h4 : _ans_10_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_187 = _ans_10_leadingZeros_T_93[3] ? 6'h3 : _ans_10_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_188 = _ans_10_leadingZeros_T_93[2] ? 6'h2 : _ans_10_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_leadingZeros_T_189 = _ans_10_leadingZeros_T_93[1] ? 6'h1 : _ans_10_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_10_leadingZeros = _ans_10_leadingZeros_T_93[0] ? 6'h0 : _ans_10_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_10_expRaw_T_1 = 6'h1f - ans_10_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_10_expRaw = ans_10_isZero ? 6'h0 : _ans_10_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_10_shiftAmt_T_2 = ans_10_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_10_shiftAmt = ans_10_expRaw > 6'h3 ? _ans_10_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_10_mantissaRaw_T = ans_10_absClipped >> ans_10_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_10_mantissaRaw = _ans_10_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_10_mantissa = ans_10_expRaw >= 6'h3 ? ans_10_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_10_expAdjusted = ans_10_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_10_exp_T_4 = ans_10_expAdjusted > 7'hf ? 4'hf : ans_10_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_10_exp = ans_10_isZero ? 4'h0 : _ans_10_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_10_fp8 = {ans_10_clippedX[31],ans_10_exp,ans_10_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_11 = {24'h0,linear_bias_11}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_11 = tempSum_11 + biasExtended_11; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_11_sign = sum32_11[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_11_absX_T = ~sum32_11; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_11_absX_T_2 = _ans_11_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_11_absX = ans_11_sign ? _ans_11_absX_T_2 : sum32_11; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_11_shiftedX_T_1 = _GEN_14432 - ans_11_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_11_shiftedX_T_3 = ans_11_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_11_shiftedX = ans_11_sign ? _ans_11_shiftedX_T_1 : _ans_11_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_11_scaledX_T_1 = ans_11_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_11_scaledX = _ans_11_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_11_clippedX_T_2 = ans_11_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_11_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_11_clippedX = ans_11_scaledX > 49'h1c0 ? 49'h1c0 : _ans_11_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_11_absClipped_T_1 = ~ans_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_11_absClipped_T_3 = _ans_11_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_11_absClipped = ans_11_clippedX[31] ? _ans_11_absClipped_T_3 : ans_11_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_11_isZero = ans_11_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39835 = {{16'd0}, ans_11_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_4 = _GEN_39835 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_6 = {ans_11_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_8 = _ans_11_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_9 = _ans_11_leadingZeros_T_4 | _ans_11_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39836 = {{8'd0}, _ans_11_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_14 = _GEN_39836 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_16 = {_ans_11_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_18 = _ans_11_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_19 = _ans_11_leadingZeros_T_14 | _ans_11_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39837 = {{4'd0}, _ans_11_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_24 = _GEN_39837 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_26 = {_ans_11_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_28 = _ans_11_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_29 = _ans_11_leadingZeros_T_24 | _ans_11_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39838 = {{2'd0}, _ans_11_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_34 = _GEN_39838 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_36 = {_ans_11_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_38 = _ans_11_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_39 = _ans_11_leadingZeros_T_34 | _ans_11_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39839 = {{1'd0}, _ans_11_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_44 = _GEN_39839 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_46 = {_ans_11_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_48 = _ans_11_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_11_leadingZeros_T_49 = _ans_11_leadingZeros_T_44 | _ans_11_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39840 = {{8'd0}, ans_11_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_55 = _GEN_39840 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_57 = {ans_11_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_59 = _ans_11_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_60 = _ans_11_leadingZeros_T_55 | _ans_11_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39841 = {{4'd0}, _ans_11_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_65 = _GEN_39841 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_67 = {_ans_11_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_69 = _ans_11_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_70 = _ans_11_leadingZeros_T_65 | _ans_11_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39842 = {{2'd0}, _ans_11_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_75 = _GEN_39842 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_77 = {_ans_11_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_79 = _ans_11_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_80 = _ans_11_leadingZeros_T_75 | _ans_11_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39843 = {{1'd0}, _ans_11_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_85 = _GEN_39843 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_87 = {_ans_11_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_89 = _ans_11_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_11_leadingZeros_T_90 = _ans_11_leadingZeros_T_85 | _ans_11_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_11_leadingZeros_T_93 = {_ans_11_leadingZeros_T_49,_ans_11_leadingZeros_T_90,ans_11_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_11_leadingZeros_T_143 = _ans_11_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_144 = _ans_11_leadingZeros_T_93[46] ? 6'h2e : _ans_11_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_145 = _ans_11_leadingZeros_T_93[45] ? 6'h2d : _ans_11_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_146 = _ans_11_leadingZeros_T_93[44] ? 6'h2c : _ans_11_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_147 = _ans_11_leadingZeros_T_93[43] ? 6'h2b : _ans_11_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_148 = _ans_11_leadingZeros_T_93[42] ? 6'h2a : _ans_11_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_149 = _ans_11_leadingZeros_T_93[41] ? 6'h29 : _ans_11_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_150 = _ans_11_leadingZeros_T_93[40] ? 6'h28 : _ans_11_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_151 = _ans_11_leadingZeros_T_93[39] ? 6'h27 : _ans_11_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_152 = _ans_11_leadingZeros_T_93[38] ? 6'h26 : _ans_11_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_153 = _ans_11_leadingZeros_T_93[37] ? 6'h25 : _ans_11_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_154 = _ans_11_leadingZeros_T_93[36] ? 6'h24 : _ans_11_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_155 = _ans_11_leadingZeros_T_93[35] ? 6'h23 : _ans_11_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_156 = _ans_11_leadingZeros_T_93[34] ? 6'h22 : _ans_11_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_157 = _ans_11_leadingZeros_T_93[33] ? 6'h21 : _ans_11_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_158 = _ans_11_leadingZeros_T_93[32] ? 6'h20 : _ans_11_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_159 = _ans_11_leadingZeros_T_93[31] ? 6'h1f : _ans_11_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_160 = _ans_11_leadingZeros_T_93[30] ? 6'h1e : _ans_11_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_161 = _ans_11_leadingZeros_T_93[29] ? 6'h1d : _ans_11_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_162 = _ans_11_leadingZeros_T_93[28] ? 6'h1c : _ans_11_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_163 = _ans_11_leadingZeros_T_93[27] ? 6'h1b : _ans_11_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_164 = _ans_11_leadingZeros_T_93[26] ? 6'h1a : _ans_11_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_165 = _ans_11_leadingZeros_T_93[25] ? 6'h19 : _ans_11_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_166 = _ans_11_leadingZeros_T_93[24] ? 6'h18 : _ans_11_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_167 = _ans_11_leadingZeros_T_93[23] ? 6'h17 : _ans_11_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_168 = _ans_11_leadingZeros_T_93[22] ? 6'h16 : _ans_11_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_169 = _ans_11_leadingZeros_T_93[21] ? 6'h15 : _ans_11_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_170 = _ans_11_leadingZeros_T_93[20] ? 6'h14 : _ans_11_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_171 = _ans_11_leadingZeros_T_93[19] ? 6'h13 : _ans_11_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_172 = _ans_11_leadingZeros_T_93[18] ? 6'h12 : _ans_11_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_173 = _ans_11_leadingZeros_T_93[17] ? 6'h11 : _ans_11_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_174 = _ans_11_leadingZeros_T_93[16] ? 6'h10 : _ans_11_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_175 = _ans_11_leadingZeros_T_93[15] ? 6'hf : _ans_11_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_176 = _ans_11_leadingZeros_T_93[14] ? 6'he : _ans_11_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_177 = _ans_11_leadingZeros_T_93[13] ? 6'hd : _ans_11_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_178 = _ans_11_leadingZeros_T_93[12] ? 6'hc : _ans_11_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_179 = _ans_11_leadingZeros_T_93[11] ? 6'hb : _ans_11_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_180 = _ans_11_leadingZeros_T_93[10] ? 6'ha : _ans_11_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_181 = _ans_11_leadingZeros_T_93[9] ? 6'h9 : _ans_11_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_182 = _ans_11_leadingZeros_T_93[8] ? 6'h8 : _ans_11_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_183 = _ans_11_leadingZeros_T_93[7] ? 6'h7 : _ans_11_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_184 = _ans_11_leadingZeros_T_93[6] ? 6'h6 : _ans_11_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_185 = _ans_11_leadingZeros_T_93[5] ? 6'h5 : _ans_11_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_186 = _ans_11_leadingZeros_T_93[4] ? 6'h4 : _ans_11_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_187 = _ans_11_leadingZeros_T_93[3] ? 6'h3 : _ans_11_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_188 = _ans_11_leadingZeros_T_93[2] ? 6'h2 : _ans_11_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_leadingZeros_T_189 = _ans_11_leadingZeros_T_93[1] ? 6'h1 : _ans_11_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_11_leadingZeros = _ans_11_leadingZeros_T_93[0] ? 6'h0 : _ans_11_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_11_expRaw_T_1 = 6'h1f - ans_11_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_11_expRaw = ans_11_isZero ? 6'h0 : _ans_11_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_11_shiftAmt_T_2 = ans_11_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_11_shiftAmt = ans_11_expRaw > 6'h3 ? _ans_11_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_11_mantissaRaw_T = ans_11_absClipped >> ans_11_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_11_mantissaRaw = _ans_11_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_11_mantissa = ans_11_expRaw >= 6'h3 ? ans_11_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_11_expAdjusted = ans_11_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_11_exp_T_4 = ans_11_expAdjusted > 7'hf ? 4'hf : ans_11_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_11_exp = ans_11_isZero ? 4'h0 : _ans_11_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_11_fp8 = {ans_11_clippedX[31],ans_11_exp,ans_11_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_12 = {24'h0,linear_bias_12}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_12 = tempSum_12 + biasExtended_12; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_12_sign = sum32_12[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_12_absX_T = ~sum32_12; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_12_absX_T_2 = _ans_12_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_12_absX = ans_12_sign ? _ans_12_absX_T_2 : sum32_12; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_12_shiftedX_T_1 = _GEN_14432 - ans_12_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_12_shiftedX_T_3 = ans_12_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_12_shiftedX = ans_12_sign ? _ans_12_shiftedX_T_1 : _ans_12_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_12_scaledX_T_1 = ans_12_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_12_scaledX = _ans_12_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_12_clippedX_T_2 = ans_12_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_12_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_12_clippedX = ans_12_scaledX > 49'h1c0 ? 49'h1c0 : _ans_12_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_12_absClipped_T_1 = ~ans_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_12_absClipped_T_3 = _ans_12_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_12_absClipped = ans_12_clippedX[31] ? _ans_12_absClipped_T_3 : ans_12_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_12_isZero = ans_12_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39846 = {{16'd0}, ans_12_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_4 = _GEN_39846 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_6 = {ans_12_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_8 = _ans_12_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_9 = _ans_12_leadingZeros_T_4 | _ans_12_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39847 = {{8'd0}, _ans_12_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_14 = _GEN_39847 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_16 = {_ans_12_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_18 = _ans_12_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_19 = _ans_12_leadingZeros_T_14 | _ans_12_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39848 = {{4'd0}, _ans_12_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_24 = _GEN_39848 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_26 = {_ans_12_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_28 = _ans_12_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_29 = _ans_12_leadingZeros_T_24 | _ans_12_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39849 = {{2'd0}, _ans_12_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_34 = _GEN_39849 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_36 = {_ans_12_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_38 = _ans_12_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_39 = _ans_12_leadingZeros_T_34 | _ans_12_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39850 = {{1'd0}, _ans_12_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_44 = _GEN_39850 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_46 = {_ans_12_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_48 = _ans_12_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_12_leadingZeros_T_49 = _ans_12_leadingZeros_T_44 | _ans_12_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39851 = {{8'd0}, ans_12_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_55 = _GEN_39851 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_57 = {ans_12_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_59 = _ans_12_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_60 = _ans_12_leadingZeros_T_55 | _ans_12_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39852 = {{4'd0}, _ans_12_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_65 = _GEN_39852 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_67 = {_ans_12_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_69 = _ans_12_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_70 = _ans_12_leadingZeros_T_65 | _ans_12_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39853 = {{2'd0}, _ans_12_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_75 = _GEN_39853 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_77 = {_ans_12_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_79 = _ans_12_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_80 = _ans_12_leadingZeros_T_75 | _ans_12_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39854 = {{1'd0}, _ans_12_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_85 = _GEN_39854 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_87 = {_ans_12_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_89 = _ans_12_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_12_leadingZeros_T_90 = _ans_12_leadingZeros_T_85 | _ans_12_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_12_leadingZeros_T_93 = {_ans_12_leadingZeros_T_49,_ans_12_leadingZeros_T_90,ans_12_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_12_leadingZeros_T_143 = _ans_12_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_144 = _ans_12_leadingZeros_T_93[46] ? 6'h2e : _ans_12_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_145 = _ans_12_leadingZeros_T_93[45] ? 6'h2d : _ans_12_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_146 = _ans_12_leadingZeros_T_93[44] ? 6'h2c : _ans_12_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_147 = _ans_12_leadingZeros_T_93[43] ? 6'h2b : _ans_12_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_148 = _ans_12_leadingZeros_T_93[42] ? 6'h2a : _ans_12_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_149 = _ans_12_leadingZeros_T_93[41] ? 6'h29 : _ans_12_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_150 = _ans_12_leadingZeros_T_93[40] ? 6'h28 : _ans_12_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_151 = _ans_12_leadingZeros_T_93[39] ? 6'h27 : _ans_12_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_152 = _ans_12_leadingZeros_T_93[38] ? 6'h26 : _ans_12_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_153 = _ans_12_leadingZeros_T_93[37] ? 6'h25 : _ans_12_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_154 = _ans_12_leadingZeros_T_93[36] ? 6'h24 : _ans_12_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_155 = _ans_12_leadingZeros_T_93[35] ? 6'h23 : _ans_12_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_156 = _ans_12_leadingZeros_T_93[34] ? 6'h22 : _ans_12_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_157 = _ans_12_leadingZeros_T_93[33] ? 6'h21 : _ans_12_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_158 = _ans_12_leadingZeros_T_93[32] ? 6'h20 : _ans_12_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_159 = _ans_12_leadingZeros_T_93[31] ? 6'h1f : _ans_12_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_160 = _ans_12_leadingZeros_T_93[30] ? 6'h1e : _ans_12_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_161 = _ans_12_leadingZeros_T_93[29] ? 6'h1d : _ans_12_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_162 = _ans_12_leadingZeros_T_93[28] ? 6'h1c : _ans_12_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_163 = _ans_12_leadingZeros_T_93[27] ? 6'h1b : _ans_12_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_164 = _ans_12_leadingZeros_T_93[26] ? 6'h1a : _ans_12_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_165 = _ans_12_leadingZeros_T_93[25] ? 6'h19 : _ans_12_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_166 = _ans_12_leadingZeros_T_93[24] ? 6'h18 : _ans_12_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_167 = _ans_12_leadingZeros_T_93[23] ? 6'h17 : _ans_12_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_168 = _ans_12_leadingZeros_T_93[22] ? 6'h16 : _ans_12_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_169 = _ans_12_leadingZeros_T_93[21] ? 6'h15 : _ans_12_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_170 = _ans_12_leadingZeros_T_93[20] ? 6'h14 : _ans_12_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_171 = _ans_12_leadingZeros_T_93[19] ? 6'h13 : _ans_12_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_172 = _ans_12_leadingZeros_T_93[18] ? 6'h12 : _ans_12_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_173 = _ans_12_leadingZeros_T_93[17] ? 6'h11 : _ans_12_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_174 = _ans_12_leadingZeros_T_93[16] ? 6'h10 : _ans_12_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_175 = _ans_12_leadingZeros_T_93[15] ? 6'hf : _ans_12_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_176 = _ans_12_leadingZeros_T_93[14] ? 6'he : _ans_12_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_177 = _ans_12_leadingZeros_T_93[13] ? 6'hd : _ans_12_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_178 = _ans_12_leadingZeros_T_93[12] ? 6'hc : _ans_12_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_179 = _ans_12_leadingZeros_T_93[11] ? 6'hb : _ans_12_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_180 = _ans_12_leadingZeros_T_93[10] ? 6'ha : _ans_12_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_181 = _ans_12_leadingZeros_T_93[9] ? 6'h9 : _ans_12_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_182 = _ans_12_leadingZeros_T_93[8] ? 6'h8 : _ans_12_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_183 = _ans_12_leadingZeros_T_93[7] ? 6'h7 : _ans_12_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_184 = _ans_12_leadingZeros_T_93[6] ? 6'h6 : _ans_12_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_185 = _ans_12_leadingZeros_T_93[5] ? 6'h5 : _ans_12_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_186 = _ans_12_leadingZeros_T_93[4] ? 6'h4 : _ans_12_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_187 = _ans_12_leadingZeros_T_93[3] ? 6'h3 : _ans_12_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_188 = _ans_12_leadingZeros_T_93[2] ? 6'h2 : _ans_12_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_leadingZeros_T_189 = _ans_12_leadingZeros_T_93[1] ? 6'h1 : _ans_12_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_12_leadingZeros = _ans_12_leadingZeros_T_93[0] ? 6'h0 : _ans_12_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_12_expRaw_T_1 = 6'h1f - ans_12_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_12_expRaw = ans_12_isZero ? 6'h0 : _ans_12_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_12_shiftAmt_T_2 = ans_12_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_12_shiftAmt = ans_12_expRaw > 6'h3 ? _ans_12_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_12_mantissaRaw_T = ans_12_absClipped >> ans_12_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_12_mantissaRaw = _ans_12_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_12_mantissa = ans_12_expRaw >= 6'h3 ? ans_12_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_12_expAdjusted = ans_12_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_12_exp_T_4 = ans_12_expAdjusted > 7'hf ? 4'hf : ans_12_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_12_exp = ans_12_isZero ? 4'h0 : _ans_12_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_12_fp8 = {ans_12_clippedX[31],ans_12_exp,ans_12_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_13 = {24'h0,linear_bias_13}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_13 = tempSum_13 + biasExtended_13; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_13_sign = sum32_13[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_13_absX_T = ~sum32_13; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_13_absX_T_2 = _ans_13_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_13_absX = ans_13_sign ? _ans_13_absX_T_2 : sum32_13; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_13_shiftedX_T_1 = _GEN_14432 - ans_13_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_13_shiftedX_T_3 = ans_13_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_13_shiftedX = ans_13_sign ? _ans_13_shiftedX_T_1 : _ans_13_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_13_scaledX_T_1 = ans_13_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_13_scaledX = _ans_13_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_13_clippedX_T_2 = ans_13_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_13_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_13_clippedX = ans_13_scaledX > 49'h1c0 ? 49'h1c0 : _ans_13_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_13_absClipped_T_1 = ~ans_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_13_absClipped_T_3 = _ans_13_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_13_absClipped = ans_13_clippedX[31] ? _ans_13_absClipped_T_3 : ans_13_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_13_isZero = ans_13_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39857 = {{16'd0}, ans_13_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_4 = _GEN_39857 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_6 = {ans_13_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_8 = _ans_13_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_9 = _ans_13_leadingZeros_T_4 | _ans_13_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39858 = {{8'd0}, _ans_13_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_14 = _GEN_39858 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_16 = {_ans_13_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_18 = _ans_13_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_19 = _ans_13_leadingZeros_T_14 | _ans_13_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39859 = {{4'd0}, _ans_13_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_24 = _GEN_39859 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_26 = {_ans_13_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_28 = _ans_13_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_29 = _ans_13_leadingZeros_T_24 | _ans_13_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39860 = {{2'd0}, _ans_13_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_34 = _GEN_39860 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_36 = {_ans_13_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_38 = _ans_13_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_39 = _ans_13_leadingZeros_T_34 | _ans_13_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39861 = {{1'd0}, _ans_13_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_44 = _GEN_39861 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_46 = {_ans_13_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_48 = _ans_13_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_13_leadingZeros_T_49 = _ans_13_leadingZeros_T_44 | _ans_13_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39862 = {{8'd0}, ans_13_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_55 = _GEN_39862 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_57 = {ans_13_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_59 = _ans_13_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_60 = _ans_13_leadingZeros_T_55 | _ans_13_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39863 = {{4'd0}, _ans_13_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_65 = _GEN_39863 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_67 = {_ans_13_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_69 = _ans_13_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_70 = _ans_13_leadingZeros_T_65 | _ans_13_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39864 = {{2'd0}, _ans_13_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_75 = _GEN_39864 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_77 = {_ans_13_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_79 = _ans_13_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_80 = _ans_13_leadingZeros_T_75 | _ans_13_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39865 = {{1'd0}, _ans_13_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_85 = _GEN_39865 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_87 = {_ans_13_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_89 = _ans_13_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_13_leadingZeros_T_90 = _ans_13_leadingZeros_T_85 | _ans_13_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_13_leadingZeros_T_93 = {_ans_13_leadingZeros_T_49,_ans_13_leadingZeros_T_90,ans_13_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_13_leadingZeros_T_143 = _ans_13_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_144 = _ans_13_leadingZeros_T_93[46] ? 6'h2e : _ans_13_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_145 = _ans_13_leadingZeros_T_93[45] ? 6'h2d : _ans_13_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_146 = _ans_13_leadingZeros_T_93[44] ? 6'h2c : _ans_13_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_147 = _ans_13_leadingZeros_T_93[43] ? 6'h2b : _ans_13_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_148 = _ans_13_leadingZeros_T_93[42] ? 6'h2a : _ans_13_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_149 = _ans_13_leadingZeros_T_93[41] ? 6'h29 : _ans_13_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_150 = _ans_13_leadingZeros_T_93[40] ? 6'h28 : _ans_13_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_151 = _ans_13_leadingZeros_T_93[39] ? 6'h27 : _ans_13_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_152 = _ans_13_leadingZeros_T_93[38] ? 6'h26 : _ans_13_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_153 = _ans_13_leadingZeros_T_93[37] ? 6'h25 : _ans_13_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_154 = _ans_13_leadingZeros_T_93[36] ? 6'h24 : _ans_13_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_155 = _ans_13_leadingZeros_T_93[35] ? 6'h23 : _ans_13_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_156 = _ans_13_leadingZeros_T_93[34] ? 6'h22 : _ans_13_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_157 = _ans_13_leadingZeros_T_93[33] ? 6'h21 : _ans_13_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_158 = _ans_13_leadingZeros_T_93[32] ? 6'h20 : _ans_13_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_159 = _ans_13_leadingZeros_T_93[31] ? 6'h1f : _ans_13_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_160 = _ans_13_leadingZeros_T_93[30] ? 6'h1e : _ans_13_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_161 = _ans_13_leadingZeros_T_93[29] ? 6'h1d : _ans_13_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_162 = _ans_13_leadingZeros_T_93[28] ? 6'h1c : _ans_13_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_163 = _ans_13_leadingZeros_T_93[27] ? 6'h1b : _ans_13_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_164 = _ans_13_leadingZeros_T_93[26] ? 6'h1a : _ans_13_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_165 = _ans_13_leadingZeros_T_93[25] ? 6'h19 : _ans_13_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_166 = _ans_13_leadingZeros_T_93[24] ? 6'h18 : _ans_13_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_167 = _ans_13_leadingZeros_T_93[23] ? 6'h17 : _ans_13_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_168 = _ans_13_leadingZeros_T_93[22] ? 6'h16 : _ans_13_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_169 = _ans_13_leadingZeros_T_93[21] ? 6'h15 : _ans_13_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_170 = _ans_13_leadingZeros_T_93[20] ? 6'h14 : _ans_13_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_171 = _ans_13_leadingZeros_T_93[19] ? 6'h13 : _ans_13_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_172 = _ans_13_leadingZeros_T_93[18] ? 6'h12 : _ans_13_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_173 = _ans_13_leadingZeros_T_93[17] ? 6'h11 : _ans_13_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_174 = _ans_13_leadingZeros_T_93[16] ? 6'h10 : _ans_13_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_175 = _ans_13_leadingZeros_T_93[15] ? 6'hf : _ans_13_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_176 = _ans_13_leadingZeros_T_93[14] ? 6'he : _ans_13_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_177 = _ans_13_leadingZeros_T_93[13] ? 6'hd : _ans_13_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_178 = _ans_13_leadingZeros_T_93[12] ? 6'hc : _ans_13_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_179 = _ans_13_leadingZeros_T_93[11] ? 6'hb : _ans_13_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_180 = _ans_13_leadingZeros_T_93[10] ? 6'ha : _ans_13_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_181 = _ans_13_leadingZeros_T_93[9] ? 6'h9 : _ans_13_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_182 = _ans_13_leadingZeros_T_93[8] ? 6'h8 : _ans_13_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_183 = _ans_13_leadingZeros_T_93[7] ? 6'h7 : _ans_13_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_184 = _ans_13_leadingZeros_T_93[6] ? 6'h6 : _ans_13_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_185 = _ans_13_leadingZeros_T_93[5] ? 6'h5 : _ans_13_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_186 = _ans_13_leadingZeros_T_93[4] ? 6'h4 : _ans_13_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_187 = _ans_13_leadingZeros_T_93[3] ? 6'h3 : _ans_13_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_188 = _ans_13_leadingZeros_T_93[2] ? 6'h2 : _ans_13_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_leadingZeros_T_189 = _ans_13_leadingZeros_T_93[1] ? 6'h1 : _ans_13_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_13_leadingZeros = _ans_13_leadingZeros_T_93[0] ? 6'h0 : _ans_13_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_13_expRaw_T_1 = 6'h1f - ans_13_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_13_expRaw = ans_13_isZero ? 6'h0 : _ans_13_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_13_shiftAmt_T_2 = ans_13_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_13_shiftAmt = ans_13_expRaw > 6'h3 ? _ans_13_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_13_mantissaRaw_T = ans_13_absClipped >> ans_13_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_13_mantissaRaw = _ans_13_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_13_mantissa = ans_13_expRaw >= 6'h3 ? ans_13_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_13_expAdjusted = ans_13_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_13_exp_T_4 = ans_13_expAdjusted > 7'hf ? 4'hf : ans_13_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_13_exp = ans_13_isZero ? 4'h0 : _ans_13_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_13_fp8 = {ans_13_clippedX[31],ans_13_exp,ans_13_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_14 = {24'h0,linear_bias_14}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_14 = tempSum_14 + biasExtended_14; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_14_sign = sum32_14[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_14_absX_T = ~sum32_14; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_14_absX_T_2 = _ans_14_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_14_absX = ans_14_sign ? _ans_14_absX_T_2 : sum32_14; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_14_shiftedX_T_1 = _GEN_14432 - ans_14_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_14_shiftedX_T_3 = ans_14_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_14_shiftedX = ans_14_sign ? _ans_14_shiftedX_T_1 : _ans_14_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_14_scaledX_T_1 = ans_14_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_14_scaledX = _ans_14_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_14_clippedX_T_2 = ans_14_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_14_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_14_clippedX = ans_14_scaledX > 49'h1c0 ? 49'h1c0 : _ans_14_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_14_absClipped_T_1 = ~ans_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_14_absClipped_T_3 = _ans_14_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_14_absClipped = ans_14_clippedX[31] ? _ans_14_absClipped_T_3 : ans_14_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_14_isZero = ans_14_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39868 = {{16'd0}, ans_14_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_4 = _GEN_39868 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_6 = {ans_14_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_8 = _ans_14_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_9 = _ans_14_leadingZeros_T_4 | _ans_14_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39869 = {{8'd0}, _ans_14_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_14 = _GEN_39869 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_16 = {_ans_14_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_18 = _ans_14_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_19 = _ans_14_leadingZeros_T_14 | _ans_14_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39870 = {{4'd0}, _ans_14_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_24 = _GEN_39870 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_26 = {_ans_14_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_28 = _ans_14_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_29 = _ans_14_leadingZeros_T_24 | _ans_14_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39871 = {{2'd0}, _ans_14_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_34 = _GEN_39871 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_36 = {_ans_14_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_38 = _ans_14_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_39 = _ans_14_leadingZeros_T_34 | _ans_14_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39872 = {{1'd0}, _ans_14_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_44 = _GEN_39872 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_46 = {_ans_14_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_48 = _ans_14_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_14_leadingZeros_T_49 = _ans_14_leadingZeros_T_44 | _ans_14_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39873 = {{8'd0}, ans_14_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_55 = _GEN_39873 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_57 = {ans_14_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_59 = _ans_14_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_60 = _ans_14_leadingZeros_T_55 | _ans_14_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39874 = {{4'd0}, _ans_14_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_65 = _GEN_39874 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_67 = {_ans_14_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_69 = _ans_14_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_70 = _ans_14_leadingZeros_T_65 | _ans_14_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39875 = {{2'd0}, _ans_14_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_75 = _GEN_39875 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_77 = {_ans_14_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_79 = _ans_14_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_80 = _ans_14_leadingZeros_T_75 | _ans_14_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39876 = {{1'd0}, _ans_14_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_85 = _GEN_39876 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_87 = {_ans_14_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_89 = _ans_14_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_14_leadingZeros_T_90 = _ans_14_leadingZeros_T_85 | _ans_14_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_14_leadingZeros_T_93 = {_ans_14_leadingZeros_T_49,_ans_14_leadingZeros_T_90,ans_14_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_14_leadingZeros_T_143 = _ans_14_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_144 = _ans_14_leadingZeros_T_93[46] ? 6'h2e : _ans_14_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_145 = _ans_14_leadingZeros_T_93[45] ? 6'h2d : _ans_14_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_146 = _ans_14_leadingZeros_T_93[44] ? 6'h2c : _ans_14_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_147 = _ans_14_leadingZeros_T_93[43] ? 6'h2b : _ans_14_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_148 = _ans_14_leadingZeros_T_93[42] ? 6'h2a : _ans_14_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_149 = _ans_14_leadingZeros_T_93[41] ? 6'h29 : _ans_14_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_150 = _ans_14_leadingZeros_T_93[40] ? 6'h28 : _ans_14_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_151 = _ans_14_leadingZeros_T_93[39] ? 6'h27 : _ans_14_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_152 = _ans_14_leadingZeros_T_93[38] ? 6'h26 : _ans_14_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_153 = _ans_14_leadingZeros_T_93[37] ? 6'h25 : _ans_14_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_154 = _ans_14_leadingZeros_T_93[36] ? 6'h24 : _ans_14_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_155 = _ans_14_leadingZeros_T_93[35] ? 6'h23 : _ans_14_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_156 = _ans_14_leadingZeros_T_93[34] ? 6'h22 : _ans_14_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_157 = _ans_14_leadingZeros_T_93[33] ? 6'h21 : _ans_14_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_158 = _ans_14_leadingZeros_T_93[32] ? 6'h20 : _ans_14_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_159 = _ans_14_leadingZeros_T_93[31] ? 6'h1f : _ans_14_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_160 = _ans_14_leadingZeros_T_93[30] ? 6'h1e : _ans_14_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_161 = _ans_14_leadingZeros_T_93[29] ? 6'h1d : _ans_14_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_162 = _ans_14_leadingZeros_T_93[28] ? 6'h1c : _ans_14_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_163 = _ans_14_leadingZeros_T_93[27] ? 6'h1b : _ans_14_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_164 = _ans_14_leadingZeros_T_93[26] ? 6'h1a : _ans_14_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_165 = _ans_14_leadingZeros_T_93[25] ? 6'h19 : _ans_14_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_166 = _ans_14_leadingZeros_T_93[24] ? 6'h18 : _ans_14_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_167 = _ans_14_leadingZeros_T_93[23] ? 6'h17 : _ans_14_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_168 = _ans_14_leadingZeros_T_93[22] ? 6'h16 : _ans_14_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_169 = _ans_14_leadingZeros_T_93[21] ? 6'h15 : _ans_14_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_170 = _ans_14_leadingZeros_T_93[20] ? 6'h14 : _ans_14_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_171 = _ans_14_leadingZeros_T_93[19] ? 6'h13 : _ans_14_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_172 = _ans_14_leadingZeros_T_93[18] ? 6'h12 : _ans_14_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_173 = _ans_14_leadingZeros_T_93[17] ? 6'h11 : _ans_14_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_174 = _ans_14_leadingZeros_T_93[16] ? 6'h10 : _ans_14_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_175 = _ans_14_leadingZeros_T_93[15] ? 6'hf : _ans_14_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_176 = _ans_14_leadingZeros_T_93[14] ? 6'he : _ans_14_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_177 = _ans_14_leadingZeros_T_93[13] ? 6'hd : _ans_14_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_178 = _ans_14_leadingZeros_T_93[12] ? 6'hc : _ans_14_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_179 = _ans_14_leadingZeros_T_93[11] ? 6'hb : _ans_14_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_180 = _ans_14_leadingZeros_T_93[10] ? 6'ha : _ans_14_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_181 = _ans_14_leadingZeros_T_93[9] ? 6'h9 : _ans_14_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_182 = _ans_14_leadingZeros_T_93[8] ? 6'h8 : _ans_14_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_183 = _ans_14_leadingZeros_T_93[7] ? 6'h7 : _ans_14_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_184 = _ans_14_leadingZeros_T_93[6] ? 6'h6 : _ans_14_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_185 = _ans_14_leadingZeros_T_93[5] ? 6'h5 : _ans_14_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_186 = _ans_14_leadingZeros_T_93[4] ? 6'h4 : _ans_14_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_187 = _ans_14_leadingZeros_T_93[3] ? 6'h3 : _ans_14_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_188 = _ans_14_leadingZeros_T_93[2] ? 6'h2 : _ans_14_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_leadingZeros_T_189 = _ans_14_leadingZeros_T_93[1] ? 6'h1 : _ans_14_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_14_leadingZeros = _ans_14_leadingZeros_T_93[0] ? 6'h0 : _ans_14_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_14_expRaw_T_1 = 6'h1f - ans_14_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_14_expRaw = ans_14_isZero ? 6'h0 : _ans_14_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_14_shiftAmt_T_2 = ans_14_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_14_shiftAmt = ans_14_expRaw > 6'h3 ? _ans_14_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_14_mantissaRaw_T = ans_14_absClipped >> ans_14_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_14_mantissaRaw = _ans_14_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_14_mantissa = ans_14_expRaw >= 6'h3 ? ans_14_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_14_expAdjusted = ans_14_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_14_exp_T_4 = ans_14_expAdjusted > 7'hf ? 4'hf : ans_14_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_14_exp = ans_14_isZero ? 4'h0 : _ans_14_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_14_fp8 = {ans_14_clippedX[31],ans_14_exp,ans_14_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_15 = {24'h0,linear_bias_15}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_15 = tempSum_15 + biasExtended_15; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_15_sign = sum32_15[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_15_absX_T = ~sum32_15; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_15_absX_T_2 = _ans_15_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_15_absX = ans_15_sign ? _ans_15_absX_T_2 : sum32_15; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_15_shiftedX_T_1 = _GEN_14432 - ans_15_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_15_shiftedX_T_3 = ans_15_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_15_shiftedX = ans_15_sign ? _ans_15_shiftedX_T_1 : _ans_15_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_15_scaledX_T_1 = ans_15_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_15_scaledX = _ans_15_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_15_clippedX_T_2 = ans_15_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_15_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_15_clippedX = ans_15_scaledX > 49'h1c0 ? 49'h1c0 : _ans_15_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_15_absClipped_T_1 = ~ans_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_15_absClipped_T_3 = _ans_15_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_15_absClipped = ans_15_clippedX[31] ? _ans_15_absClipped_T_3 : ans_15_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_15_isZero = ans_15_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39879 = {{16'd0}, ans_15_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_4 = _GEN_39879 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_6 = {ans_15_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_8 = _ans_15_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_9 = _ans_15_leadingZeros_T_4 | _ans_15_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39880 = {{8'd0}, _ans_15_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_14 = _GEN_39880 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_16 = {_ans_15_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_18 = _ans_15_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_19 = _ans_15_leadingZeros_T_14 | _ans_15_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39881 = {{4'd0}, _ans_15_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_24 = _GEN_39881 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_26 = {_ans_15_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_28 = _ans_15_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_29 = _ans_15_leadingZeros_T_24 | _ans_15_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39882 = {{2'd0}, _ans_15_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_34 = _GEN_39882 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_36 = {_ans_15_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_38 = _ans_15_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_39 = _ans_15_leadingZeros_T_34 | _ans_15_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39883 = {{1'd0}, _ans_15_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_44 = _GEN_39883 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_46 = {_ans_15_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_48 = _ans_15_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_15_leadingZeros_T_49 = _ans_15_leadingZeros_T_44 | _ans_15_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39884 = {{8'd0}, ans_15_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_55 = _GEN_39884 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_57 = {ans_15_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_59 = _ans_15_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_60 = _ans_15_leadingZeros_T_55 | _ans_15_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39885 = {{4'd0}, _ans_15_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_65 = _GEN_39885 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_67 = {_ans_15_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_69 = _ans_15_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_70 = _ans_15_leadingZeros_T_65 | _ans_15_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39886 = {{2'd0}, _ans_15_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_75 = _GEN_39886 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_77 = {_ans_15_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_79 = _ans_15_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_80 = _ans_15_leadingZeros_T_75 | _ans_15_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39887 = {{1'd0}, _ans_15_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_85 = _GEN_39887 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_87 = {_ans_15_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_89 = _ans_15_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_15_leadingZeros_T_90 = _ans_15_leadingZeros_T_85 | _ans_15_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_15_leadingZeros_T_93 = {_ans_15_leadingZeros_T_49,_ans_15_leadingZeros_T_90,ans_15_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_15_leadingZeros_T_143 = _ans_15_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_144 = _ans_15_leadingZeros_T_93[46] ? 6'h2e : _ans_15_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_145 = _ans_15_leadingZeros_T_93[45] ? 6'h2d : _ans_15_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_146 = _ans_15_leadingZeros_T_93[44] ? 6'h2c : _ans_15_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_147 = _ans_15_leadingZeros_T_93[43] ? 6'h2b : _ans_15_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_148 = _ans_15_leadingZeros_T_93[42] ? 6'h2a : _ans_15_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_149 = _ans_15_leadingZeros_T_93[41] ? 6'h29 : _ans_15_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_150 = _ans_15_leadingZeros_T_93[40] ? 6'h28 : _ans_15_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_151 = _ans_15_leadingZeros_T_93[39] ? 6'h27 : _ans_15_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_152 = _ans_15_leadingZeros_T_93[38] ? 6'h26 : _ans_15_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_153 = _ans_15_leadingZeros_T_93[37] ? 6'h25 : _ans_15_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_154 = _ans_15_leadingZeros_T_93[36] ? 6'h24 : _ans_15_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_155 = _ans_15_leadingZeros_T_93[35] ? 6'h23 : _ans_15_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_156 = _ans_15_leadingZeros_T_93[34] ? 6'h22 : _ans_15_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_157 = _ans_15_leadingZeros_T_93[33] ? 6'h21 : _ans_15_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_158 = _ans_15_leadingZeros_T_93[32] ? 6'h20 : _ans_15_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_159 = _ans_15_leadingZeros_T_93[31] ? 6'h1f : _ans_15_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_160 = _ans_15_leadingZeros_T_93[30] ? 6'h1e : _ans_15_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_161 = _ans_15_leadingZeros_T_93[29] ? 6'h1d : _ans_15_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_162 = _ans_15_leadingZeros_T_93[28] ? 6'h1c : _ans_15_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_163 = _ans_15_leadingZeros_T_93[27] ? 6'h1b : _ans_15_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_164 = _ans_15_leadingZeros_T_93[26] ? 6'h1a : _ans_15_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_165 = _ans_15_leadingZeros_T_93[25] ? 6'h19 : _ans_15_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_166 = _ans_15_leadingZeros_T_93[24] ? 6'h18 : _ans_15_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_167 = _ans_15_leadingZeros_T_93[23] ? 6'h17 : _ans_15_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_168 = _ans_15_leadingZeros_T_93[22] ? 6'h16 : _ans_15_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_169 = _ans_15_leadingZeros_T_93[21] ? 6'h15 : _ans_15_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_170 = _ans_15_leadingZeros_T_93[20] ? 6'h14 : _ans_15_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_171 = _ans_15_leadingZeros_T_93[19] ? 6'h13 : _ans_15_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_172 = _ans_15_leadingZeros_T_93[18] ? 6'h12 : _ans_15_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_173 = _ans_15_leadingZeros_T_93[17] ? 6'h11 : _ans_15_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_174 = _ans_15_leadingZeros_T_93[16] ? 6'h10 : _ans_15_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_175 = _ans_15_leadingZeros_T_93[15] ? 6'hf : _ans_15_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_176 = _ans_15_leadingZeros_T_93[14] ? 6'he : _ans_15_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_177 = _ans_15_leadingZeros_T_93[13] ? 6'hd : _ans_15_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_178 = _ans_15_leadingZeros_T_93[12] ? 6'hc : _ans_15_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_179 = _ans_15_leadingZeros_T_93[11] ? 6'hb : _ans_15_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_180 = _ans_15_leadingZeros_T_93[10] ? 6'ha : _ans_15_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_181 = _ans_15_leadingZeros_T_93[9] ? 6'h9 : _ans_15_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_182 = _ans_15_leadingZeros_T_93[8] ? 6'h8 : _ans_15_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_183 = _ans_15_leadingZeros_T_93[7] ? 6'h7 : _ans_15_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_184 = _ans_15_leadingZeros_T_93[6] ? 6'h6 : _ans_15_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_185 = _ans_15_leadingZeros_T_93[5] ? 6'h5 : _ans_15_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_186 = _ans_15_leadingZeros_T_93[4] ? 6'h4 : _ans_15_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_187 = _ans_15_leadingZeros_T_93[3] ? 6'h3 : _ans_15_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_188 = _ans_15_leadingZeros_T_93[2] ? 6'h2 : _ans_15_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_leadingZeros_T_189 = _ans_15_leadingZeros_T_93[1] ? 6'h1 : _ans_15_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_15_leadingZeros = _ans_15_leadingZeros_T_93[0] ? 6'h0 : _ans_15_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_15_expRaw_T_1 = 6'h1f - ans_15_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_15_expRaw = ans_15_isZero ? 6'h0 : _ans_15_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_15_shiftAmt_T_2 = ans_15_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_15_shiftAmt = ans_15_expRaw > 6'h3 ? _ans_15_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_15_mantissaRaw_T = ans_15_absClipped >> ans_15_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_15_mantissaRaw = _ans_15_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_15_mantissa = ans_15_expRaw >= 6'h3 ? ans_15_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_15_expAdjusted = ans_15_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_15_exp_T_4 = ans_15_expAdjusted > 7'hf ? 4'hf : ans_15_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_15_exp = ans_15_isZero ? 4'h0 : _ans_15_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_15_fp8 = {ans_15_clippedX[31],ans_15_exp,ans_15_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_16 = {24'h0,linear_bias_16}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_16 = tempSum_16 + biasExtended_16; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_16_sign = sum32_16[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_16_absX_T = ~sum32_16; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_16_absX_T_2 = _ans_16_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_16_absX = ans_16_sign ? _ans_16_absX_T_2 : sum32_16; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_16_shiftedX_T_1 = _GEN_14432 - ans_16_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_16_shiftedX_T_3 = ans_16_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_16_shiftedX = ans_16_sign ? _ans_16_shiftedX_T_1 : _ans_16_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_16_scaledX_T_1 = ans_16_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_16_scaledX = _ans_16_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_16_clippedX_T_2 = ans_16_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_16_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_16_clippedX = ans_16_scaledX > 49'h1c0 ? 49'h1c0 : _ans_16_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_16_absClipped_T_1 = ~ans_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_16_absClipped_T_3 = _ans_16_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_16_absClipped = ans_16_clippedX[31] ? _ans_16_absClipped_T_3 : ans_16_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_16_isZero = ans_16_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39890 = {{16'd0}, ans_16_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_4 = _GEN_39890 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_6 = {ans_16_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_8 = _ans_16_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_9 = _ans_16_leadingZeros_T_4 | _ans_16_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39891 = {{8'd0}, _ans_16_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_14 = _GEN_39891 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_16 = {_ans_16_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_18 = _ans_16_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_19 = _ans_16_leadingZeros_T_14 | _ans_16_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39892 = {{4'd0}, _ans_16_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_24 = _GEN_39892 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_26 = {_ans_16_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_28 = _ans_16_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_29 = _ans_16_leadingZeros_T_24 | _ans_16_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39893 = {{2'd0}, _ans_16_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_34 = _GEN_39893 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_36 = {_ans_16_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_38 = _ans_16_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_39 = _ans_16_leadingZeros_T_34 | _ans_16_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39894 = {{1'd0}, _ans_16_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_44 = _GEN_39894 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_46 = {_ans_16_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_48 = _ans_16_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_16_leadingZeros_T_49 = _ans_16_leadingZeros_T_44 | _ans_16_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39895 = {{8'd0}, ans_16_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_55 = _GEN_39895 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_57 = {ans_16_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_59 = _ans_16_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_60 = _ans_16_leadingZeros_T_55 | _ans_16_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39896 = {{4'd0}, _ans_16_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_65 = _GEN_39896 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_67 = {_ans_16_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_69 = _ans_16_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_70 = _ans_16_leadingZeros_T_65 | _ans_16_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39897 = {{2'd0}, _ans_16_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_75 = _GEN_39897 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_77 = {_ans_16_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_79 = _ans_16_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_80 = _ans_16_leadingZeros_T_75 | _ans_16_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39898 = {{1'd0}, _ans_16_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_85 = _GEN_39898 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_87 = {_ans_16_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_89 = _ans_16_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_16_leadingZeros_T_90 = _ans_16_leadingZeros_T_85 | _ans_16_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_16_leadingZeros_T_93 = {_ans_16_leadingZeros_T_49,_ans_16_leadingZeros_T_90,ans_16_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_16_leadingZeros_T_143 = _ans_16_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_144 = _ans_16_leadingZeros_T_93[46] ? 6'h2e : _ans_16_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_145 = _ans_16_leadingZeros_T_93[45] ? 6'h2d : _ans_16_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_146 = _ans_16_leadingZeros_T_93[44] ? 6'h2c : _ans_16_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_147 = _ans_16_leadingZeros_T_93[43] ? 6'h2b : _ans_16_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_148 = _ans_16_leadingZeros_T_93[42] ? 6'h2a : _ans_16_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_149 = _ans_16_leadingZeros_T_93[41] ? 6'h29 : _ans_16_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_150 = _ans_16_leadingZeros_T_93[40] ? 6'h28 : _ans_16_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_151 = _ans_16_leadingZeros_T_93[39] ? 6'h27 : _ans_16_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_152 = _ans_16_leadingZeros_T_93[38] ? 6'h26 : _ans_16_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_153 = _ans_16_leadingZeros_T_93[37] ? 6'h25 : _ans_16_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_154 = _ans_16_leadingZeros_T_93[36] ? 6'h24 : _ans_16_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_155 = _ans_16_leadingZeros_T_93[35] ? 6'h23 : _ans_16_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_156 = _ans_16_leadingZeros_T_93[34] ? 6'h22 : _ans_16_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_157 = _ans_16_leadingZeros_T_93[33] ? 6'h21 : _ans_16_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_158 = _ans_16_leadingZeros_T_93[32] ? 6'h20 : _ans_16_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_159 = _ans_16_leadingZeros_T_93[31] ? 6'h1f : _ans_16_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_160 = _ans_16_leadingZeros_T_93[30] ? 6'h1e : _ans_16_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_161 = _ans_16_leadingZeros_T_93[29] ? 6'h1d : _ans_16_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_162 = _ans_16_leadingZeros_T_93[28] ? 6'h1c : _ans_16_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_163 = _ans_16_leadingZeros_T_93[27] ? 6'h1b : _ans_16_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_164 = _ans_16_leadingZeros_T_93[26] ? 6'h1a : _ans_16_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_165 = _ans_16_leadingZeros_T_93[25] ? 6'h19 : _ans_16_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_166 = _ans_16_leadingZeros_T_93[24] ? 6'h18 : _ans_16_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_167 = _ans_16_leadingZeros_T_93[23] ? 6'h17 : _ans_16_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_168 = _ans_16_leadingZeros_T_93[22] ? 6'h16 : _ans_16_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_169 = _ans_16_leadingZeros_T_93[21] ? 6'h15 : _ans_16_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_170 = _ans_16_leadingZeros_T_93[20] ? 6'h14 : _ans_16_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_171 = _ans_16_leadingZeros_T_93[19] ? 6'h13 : _ans_16_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_172 = _ans_16_leadingZeros_T_93[18] ? 6'h12 : _ans_16_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_173 = _ans_16_leadingZeros_T_93[17] ? 6'h11 : _ans_16_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_174 = _ans_16_leadingZeros_T_93[16] ? 6'h10 : _ans_16_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_175 = _ans_16_leadingZeros_T_93[15] ? 6'hf : _ans_16_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_176 = _ans_16_leadingZeros_T_93[14] ? 6'he : _ans_16_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_177 = _ans_16_leadingZeros_T_93[13] ? 6'hd : _ans_16_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_178 = _ans_16_leadingZeros_T_93[12] ? 6'hc : _ans_16_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_179 = _ans_16_leadingZeros_T_93[11] ? 6'hb : _ans_16_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_180 = _ans_16_leadingZeros_T_93[10] ? 6'ha : _ans_16_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_181 = _ans_16_leadingZeros_T_93[9] ? 6'h9 : _ans_16_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_182 = _ans_16_leadingZeros_T_93[8] ? 6'h8 : _ans_16_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_183 = _ans_16_leadingZeros_T_93[7] ? 6'h7 : _ans_16_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_184 = _ans_16_leadingZeros_T_93[6] ? 6'h6 : _ans_16_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_185 = _ans_16_leadingZeros_T_93[5] ? 6'h5 : _ans_16_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_186 = _ans_16_leadingZeros_T_93[4] ? 6'h4 : _ans_16_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_187 = _ans_16_leadingZeros_T_93[3] ? 6'h3 : _ans_16_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_188 = _ans_16_leadingZeros_T_93[2] ? 6'h2 : _ans_16_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_leadingZeros_T_189 = _ans_16_leadingZeros_T_93[1] ? 6'h1 : _ans_16_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_16_leadingZeros = _ans_16_leadingZeros_T_93[0] ? 6'h0 : _ans_16_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_16_expRaw_T_1 = 6'h1f - ans_16_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_16_expRaw = ans_16_isZero ? 6'h0 : _ans_16_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_16_shiftAmt_T_2 = ans_16_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_16_shiftAmt = ans_16_expRaw > 6'h3 ? _ans_16_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_16_mantissaRaw_T = ans_16_absClipped >> ans_16_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_16_mantissaRaw = _ans_16_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_16_mantissa = ans_16_expRaw >= 6'h3 ? ans_16_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_16_expAdjusted = ans_16_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_16_exp_T_4 = ans_16_expAdjusted > 7'hf ? 4'hf : ans_16_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_16_exp = ans_16_isZero ? 4'h0 : _ans_16_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_16_fp8 = {ans_16_clippedX[31],ans_16_exp,ans_16_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_17 = {24'h0,linear_bias_17}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_17 = tempSum_17 + biasExtended_17; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_17_sign = sum32_17[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_17_absX_T = ~sum32_17; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_17_absX_T_2 = _ans_17_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_17_absX = ans_17_sign ? _ans_17_absX_T_2 : sum32_17; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_17_shiftedX_T_1 = _GEN_14432 - ans_17_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_17_shiftedX_T_3 = ans_17_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_17_shiftedX = ans_17_sign ? _ans_17_shiftedX_T_1 : _ans_17_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_17_scaledX_T_1 = ans_17_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_17_scaledX = _ans_17_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_17_clippedX_T_2 = ans_17_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_17_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_17_clippedX = ans_17_scaledX > 49'h1c0 ? 49'h1c0 : _ans_17_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_17_absClipped_T_1 = ~ans_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_17_absClipped_T_3 = _ans_17_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_17_absClipped = ans_17_clippedX[31] ? _ans_17_absClipped_T_3 : ans_17_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_17_isZero = ans_17_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39901 = {{16'd0}, ans_17_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_4 = _GEN_39901 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_6 = {ans_17_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_8 = _ans_17_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_9 = _ans_17_leadingZeros_T_4 | _ans_17_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39902 = {{8'd0}, _ans_17_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_14 = _GEN_39902 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_16 = {_ans_17_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_18 = _ans_17_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_19 = _ans_17_leadingZeros_T_14 | _ans_17_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39903 = {{4'd0}, _ans_17_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_24 = _GEN_39903 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_26 = {_ans_17_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_28 = _ans_17_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_29 = _ans_17_leadingZeros_T_24 | _ans_17_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39904 = {{2'd0}, _ans_17_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_34 = _GEN_39904 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_36 = {_ans_17_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_38 = _ans_17_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_39 = _ans_17_leadingZeros_T_34 | _ans_17_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39905 = {{1'd0}, _ans_17_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_44 = _GEN_39905 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_46 = {_ans_17_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_48 = _ans_17_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_17_leadingZeros_T_49 = _ans_17_leadingZeros_T_44 | _ans_17_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39906 = {{8'd0}, ans_17_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_55 = _GEN_39906 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_57 = {ans_17_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_59 = _ans_17_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_60 = _ans_17_leadingZeros_T_55 | _ans_17_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39907 = {{4'd0}, _ans_17_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_65 = _GEN_39907 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_67 = {_ans_17_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_69 = _ans_17_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_70 = _ans_17_leadingZeros_T_65 | _ans_17_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39908 = {{2'd0}, _ans_17_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_75 = _GEN_39908 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_77 = {_ans_17_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_79 = _ans_17_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_80 = _ans_17_leadingZeros_T_75 | _ans_17_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39909 = {{1'd0}, _ans_17_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_85 = _GEN_39909 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_87 = {_ans_17_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_89 = _ans_17_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_17_leadingZeros_T_90 = _ans_17_leadingZeros_T_85 | _ans_17_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_17_leadingZeros_T_93 = {_ans_17_leadingZeros_T_49,_ans_17_leadingZeros_T_90,ans_17_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_17_leadingZeros_T_143 = _ans_17_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_144 = _ans_17_leadingZeros_T_93[46] ? 6'h2e : _ans_17_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_145 = _ans_17_leadingZeros_T_93[45] ? 6'h2d : _ans_17_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_146 = _ans_17_leadingZeros_T_93[44] ? 6'h2c : _ans_17_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_147 = _ans_17_leadingZeros_T_93[43] ? 6'h2b : _ans_17_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_148 = _ans_17_leadingZeros_T_93[42] ? 6'h2a : _ans_17_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_149 = _ans_17_leadingZeros_T_93[41] ? 6'h29 : _ans_17_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_150 = _ans_17_leadingZeros_T_93[40] ? 6'h28 : _ans_17_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_151 = _ans_17_leadingZeros_T_93[39] ? 6'h27 : _ans_17_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_152 = _ans_17_leadingZeros_T_93[38] ? 6'h26 : _ans_17_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_153 = _ans_17_leadingZeros_T_93[37] ? 6'h25 : _ans_17_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_154 = _ans_17_leadingZeros_T_93[36] ? 6'h24 : _ans_17_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_155 = _ans_17_leadingZeros_T_93[35] ? 6'h23 : _ans_17_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_156 = _ans_17_leadingZeros_T_93[34] ? 6'h22 : _ans_17_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_157 = _ans_17_leadingZeros_T_93[33] ? 6'h21 : _ans_17_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_158 = _ans_17_leadingZeros_T_93[32] ? 6'h20 : _ans_17_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_159 = _ans_17_leadingZeros_T_93[31] ? 6'h1f : _ans_17_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_160 = _ans_17_leadingZeros_T_93[30] ? 6'h1e : _ans_17_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_161 = _ans_17_leadingZeros_T_93[29] ? 6'h1d : _ans_17_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_162 = _ans_17_leadingZeros_T_93[28] ? 6'h1c : _ans_17_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_163 = _ans_17_leadingZeros_T_93[27] ? 6'h1b : _ans_17_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_164 = _ans_17_leadingZeros_T_93[26] ? 6'h1a : _ans_17_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_165 = _ans_17_leadingZeros_T_93[25] ? 6'h19 : _ans_17_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_166 = _ans_17_leadingZeros_T_93[24] ? 6'h18 : _ans_17_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_167 = _ans_17_leadingZeros_T_93[23] ? 6'h17 : _ans_17_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_168 = _ans_17_leadingZeros_T_93[22] ? 6'h16 : _ans_17_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_169 = _ans_17_leadingZeros_T_93[21] ? 6'h15 : _ans_17_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_170 = _ans_17_leadingZeros_T_93[20] ? 6'h14 : _ans_17_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_171 = _ans_17_leadingZeros_T_93[19] ? 6'h13 : _ans_17_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_172 = _ans_17_leadingZeros_T_93[18] ? 6'h12 : _ans_17_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_173 = _ans_17_leadingZeros_T_93[17] ? 6'h11 : _ans_17_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_174 = _ans_17_leadingZeros_T_93[16] ? 6'h10 : _ans_17_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_175 = _ans_17_leadingZeros_T_93[15] ? 6'hf : _ans_17_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_176 = _ans_17_leadingZeros_T_93[14] ? 6'he : _ans_17_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_177 = _ans_17_leadingZeros_T_93[13] ? 6'hd : _ans_17_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_178 = _ans_17_leadingZeros_T_93[12] ? 6'hc : _ans_17_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_179 = _ans_17_leadingZeros_T_93[11] ? 6'hb : _ans_17_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_180 = _ans_17_leadingZeros_T_93[10] ? 6'ha : _ans_17_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_181 = _ans_17_leadingZeros_T_93[9] ? 6'h9 : _ans_17_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_182 = _ans_17_leadingZeros_T_93[8] ? 6'h8 : _ans_17_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_183 = _ans_17_leadingZeros_T_93[7] ? 6'h7 : _ans_17_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_184 = _ans_17_leadingZeros_T_93[6] ? 6'h6 : _ans_17_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_185 = _ans_17_leadingZeros_T_93[5] ? 6'h5 : _ans_17_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_186 = _ans_17_leadingZeros_T_93[4] ? 6'h4 : _ans_17_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_187 = _ans_17_leadingZeros_T_93[3] ? 6'h3 : _ans_17_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_188 = _ans_17_leadingZeros_T_93[2] ? 6'h2 : _ans_17_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_leadingZeros_T_189 = _ans_17_leadingZeros_T_93[1] ? 6'h1 : _ans_17_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_17_leadingZeros = _ans_17_leadingZeros_T_93[0] ? 6'h0 : _ans_17_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_17_expRaw_T_1 = 6'h1f - ans_17_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_17_expRaw = ans_17_isZero ? 6'h0 : _ans_17_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_17_shiftAmt_T_2 = ans_17_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_17_shiftAmt = ans_17_expRaw > 6'h3 ? _ans_17_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_17_mantissaRaw_T = ans_17_absClipped >> ans_17_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_17_mantissaRaw = _ans_17_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_17_mantissa = ans_17_expRaw >= 6'h3 ? ans_17_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_17_expAdjusted = ans_17_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_17_exp_T_4 = ans_17_expAdjusted > 7'hf ? 4'hf : ans_17_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_17_exp = ans_17_isZero ? 4'h0 : _ans_17_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_17_fp8 = {ans_17_clippedX[31],ans_17_exp,ans_17_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_18 = {24'h0,linear_bias_18}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_18 = tempSum_18 + biasExtended_18; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_18_sign = sum32_18[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_18_absX_T = ~sum32_18; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_18_absX_T_2 = _ans_18_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_18_absX = ans_18_sign ? _ans_18_absX_T_2 : sum32_18; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_18_shiftedX_T_1 = _GEN_14432 - ans_18_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_18_shiftedX_T_3 = ans_18_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_18_shiftedX = ans_18_sign ? _ans_18_shiftedX_T_1 : _ans_18_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_18_scaledX_T_1 = ans_18_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_18_scaledX = _ans_18_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_18_clippedX_T_2 = ans_18_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_18_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_18_clippedX = ans_18_scaledX > 49'h1c0 ? 49'h1c0 : _ans_18_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_18_absClipped_T_1 = ~ans_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_18_absClipped_T_3 = _ans_18_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_18_absClipped = ans_18_clippedX[31] ? _ans_18_absClipped_T_3 : ans_18_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_18_isZero = ans_18_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39912 = {{16'd0}, ans_18_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_4 = _GEN_39912 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_6 = {ans_18_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_8 = _ans_18_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_9 = _ans_18_leadingZeros_T_4 | _ans_18_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39913 = {{8'd0}, _ans_18_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_14 = _GEN_39913 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_16 = {_ans_18_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_18 = _ans_18_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_19 = _ans_18_leadingZeros_T_14 | _ans_18_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39914 = {{4'd0}, _ans_18_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_24 = _GEN_39914 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_26 = {_ans_18_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_28 = _ans_18_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_29 = _ans_18_leadingZeros_T_24 | _ans_18_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39915 = {{2'd0}, _ans_18_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_34 = _GEN_39915 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_36 = {_ans_18_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_38 = _ans_18_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_39 = _ans_18_leadingZeros_T_34 | _ans_18_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39916 = {{1'd0}, _ans_18_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_44 = _GEN_39916 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_46 = {_ans_18_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_48 = _ans_18_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_18_leadingZeros_T_49 = _ans_18_leadingZeros_T_44 | _ans_18_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39917 = {{8'd0}, ans_18_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_55 = _GEN_39917 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_57 = {ans_18_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_59 = _ans_18_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_60 = _ans_18_leadingZeros_T_55 | _ans_18_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39918 = {{4'd0}, _ans_18_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_65 = _GEN_39918 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_67 = {_ans_18_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_69 = _ans_18_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_70 = _ans_18_leadingZeros_T_65 | _ans_18_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39919 = {{2'd0}, _ans_18_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_75 = _GEN_39919 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_77 = {_ans_18_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_79 = _ans_18_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_80 = _ans_18_leadingZeros_T_75 | _ans_18_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39920 = {{1'd0}, _ans_18_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_85 = _GEN_39920 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_87 = {_ans_18_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_89 = _ans_18_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_18_leadingZeros_T_90 = _ans_18_leadingZeros_T_85 | _ans_18_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_18_leadingZeros_T_93 = {_ans_18_leadingZeros_T_49,_ans_18_leadingZeros_T_90,ans_18_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_18_leadingZeros_T_143 = _ans_18_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_144 = _ans_18_leadingZeros_T_93[46] ? 6'h2e : _ans_18_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_145 = _ans_18_leadingZeros_T_93[45] ? 6'h2d : _ans_18_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_146 = _ans_18_leadingZeros_T_93[44] ? 6'h2c : _ans_18_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_147 = _ans_18_leadingZeros_T_93[43] ? 6'h2b : _ans_18_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_148 = _ans_18_leadingZeros_T_93[42] ? 6'h2a : _ans_18_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_149 = _ans_18_leadingZeros_T_93[41] ? 6'h29 : _ans_18_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_150 = _ans_18_leadingZeros_T_93[40] ? 6'h28 : _ans_18_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_151 = _ans_18_leadingZeros_T_93[39] ? 6'h27 : _ans_18_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_152 = _ans_18_leadingZeros_T_93[38] ? 6'h26 : _ans_18_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_153 = _ans_18_leadingZeros_T_93[37] ? 6'h25 : _ans_18_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_154 = _ans_18_leadingZeros_T_93[36] ? 6'h24 : _ans_18_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_155 = _ans_18_leadingZeros_T_93[35] ? 6'h23 : _ans_18_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_156 = _ans_18_leadingZeros_T_93[34] ? 6'h22 : _ans_18_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_157 = _ans_18_leadingZeros_T_93[33] ? 6'h21 : _ans_18_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_158 = _ans_18_leadingZeros_T_93[32] ? 6'h20 : _ans_18_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_159 = _ans_18_leadingZeros_T_93[31] ? 6'h1f : _ans_18_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_160 = _ans_18_leadingZeros_T_93[30] ? 6'h1e : _ans_18_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_161 = _ans_18_leadingZeros_T_93[29] ? 6'h1d : _ans_18_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_162 = _ans_18_leadingZeros_T_93[28] ? 6'h1c : _ans_18_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_163 = _ans_18_leadingZeros_T_93[27] ? 6'h1b : _ans_18_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_164 = _ans_18_leadingZeros_T_93[26] ? 6'h1a : _ans_18_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_165 = _ans_18_leadingZeros_T_93[25] ? 6'h19 : _ans_18_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_166 = _ans_18_leadingZeros_T_93[24] ? 6'h18 : _ans_18_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_167 = _ans_18_leadingZeros_T_93[23] ? 6'h17 : _ans_18_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_168 = _ans_18_leadingZeros_T_93[22] ? 6'h16 : _ans_18_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_169 = _ans_18_leadingZeros_T_93[21] ? 6'h15 : _ans_18_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_170 = _ans_18_leadingZeros_T_93[20] ? 6'h14 : _ans_18_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_171 = _ans_18_leadingZeros_T_93[19] ? 6'h13 : _ans_18_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_172 = _ans_18_leadingZeros_T_93[18] ? 6'h12 : _ans_18_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_173 = _ans_18_leadingZeros_T_93[17] ? 6'h11 : _ans_18_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_174 = _ans_18_leadingZeros_T_93[16] ? 6'h10 : _ans_18_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_175 = _ans_18_leadingZeros_T_93[15] ? 6'hf : _ans_18_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_176 = _ans_18_leadingZeros_T_93[14] ? 6'he : _ans_18_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_177 = _ans_18_leadingZeros_T_93[13] ? 6'hd : _ans_18_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_178 = _ans_18_leadingZeros_T_93[12] ? 6'hc : _ans_18_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_179 = _ans_18_leadingZeros_T_93[11] ? 6'hb : _ans_18_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_180 = _ans_18_leadingZeros_T_93[10] ? 6'ha : _ans_18_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_181 = _ans_18_leadingZeros_T_93[9] ? 6'h9 : _ans_18_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_182 = _ans_18_leadingZeros_T_93[8] ? 6'h8 : _ans_18_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_183 = _ans_18_leadingZeros_T_93[7] ? 6'h7 : _ans_18_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_184 = _ans_18_leadingZeros_T_93[6] ? 6'h6 : _ans_18_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_185 = _ans_18_leadingZeros_T_93[5] ? 6'h5 : _ans_18_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_186 = _ans_18_leadingZeros_T_93[4] ? 6'h4 : _ans_18_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_187 = _ans_18_leadingZeros_T_93[3] ? 6'h3 : _ans_18_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_188 = _ans_18_leadingZeros_T_93[2] ? 6'h2 : _ans_18_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_leadingZeros_T_189 = _ans_18_leadingZeros_T_93[1] ? 6'h1 : _ans_18_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_18_leadingZeros = _ans_18_leadingZeros_T_93[0] ? 6'h0 : _ans_18_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_18_expRaw_T_1 = 6'h1f - ans_18_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_18_expRaw = ans_18_isZero ? 6'h0 : _ans_18_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_18_shiftAmt_T_2 = ans_18_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_18_shiftAmt = ans_18_expRaw > 6'h3 ? _ans_18_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_18_mantissaRaw_T = ans_18_absClipped >> ans_18_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_18_mantissaRaw = _ans_18_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_18_mantissa = ans_18_expRaw >= 6'h3 ? ans_18_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_18_expAdjusted = ans_18_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_18_exp_T_4 = ans_18_expAdjusted > 7'hf ? 4'hf : ans_18_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_18_exp = ans_18_isZero ? 4'h0 : _ans_18_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_18_fp8 = {ans_18_clippedX[31],ans_18_exp,ans_18_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_19 = {24'h0,linear_bias_19}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_19 = tempSum_19 + biasExtended_19; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_19_sign = sum32_19[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_19_absX_T = ~sum32_19; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_19_absX_T_2 = _ans_19_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_19_absX = ans_19_sign ? _ans_19_absX_T_2 : sum32_19; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_19_shiftedX_T_1 = _GEN_14432 - ans_19_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_19_shiftedX_T_3 = ans_19_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_19_shiftedX = ans_19_sign ? _ans_19_shiftedX_T_1 : _ans_19_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_19_scaledX_T_1 = ans_19_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_19_scaledX = _ans_19_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_19_clippedX_T_2 = ans_19_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_19_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_19_clippedX = ans_19_scaledX > 49'h1c0 ? 49'h1c0 : _ans_19_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_19_absClipped_T_1 = ~ans_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_19_absClipped_T_3 = _ans_19_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_19_absClipped = ans_19_clippedX[31] ? _ans_19_absClipped_T_3 : ans_19_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_19_isZero = ans_19_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39923 = {{16'd0}, ans_19_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_4 = _GEN_39923 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_6 = {ans_19_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_8 = _ans_19_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_9 = _ans_19_leadingZeros_T_4 | _ans_19_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39924 = {{8'd0}, _ans_19_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_14 = _GEN_39924 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_16 = {_ans_19_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_18 = _ans_19_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_19 = _ans_19_leadingZeros_T_14 | _ans_19_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39925 = {{4'd0}, _ans_19_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_24 = _GEN_39925 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_26 = {_ans_19_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_28 = _ans_19_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_29 = _ans_19_leadingZeros_T_24 | _ans_19_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39926 = {{2'd0}, _ans_19_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_34 = _GEN_39926 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_36 = {_ans_19_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_38 = _ans_19_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_39 = _ans_19_leadingZeros_T_34 | _ans_19_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39927 = {{1'd0}, _ans_19_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_44 = _GEN_39927 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_46 = {_ans_19_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_48 = _ans_19_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_19_leadingZeros_T_49 = _ans_19_leadingZeros_T_44 | _ans_19_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39928 = {{8'd0}, ans_19_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_55 = _GEN_39928 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_57 = {ans_19_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_59 = _ans_19_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_60 = _ans_19_leadingZeros_T_55 | _ans_19_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39929 = {{4'd0}, _ans_19_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_65 = _GEN_39929 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_67 = {_ans_19_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_69 = _ans_19_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_70 = _ans_19_leadingZeros_T_65 | _ans_19_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39930 = {{2'd0}, _ans_19_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_75 = _GEN_39930 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_77 = {_ans_19_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_79 = _ans_19_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_80 = _ans_19_leadingZeros_T_75 | _ans_19_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39931 = {{1'd0}, _ans_19_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_85 = _GEN_39931 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_87 = {_ans_19_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_89 = _ans_19_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_19_leadingZeros_T_90 = _ans_19_leadingZeros_T_85 | _ans_19_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_19_leadingZeros_T_93 = {_ans_19_leadingZeros_T_49,_ans_19_leadingZeros_T_90,ans_19_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_19_leadingZeros_T_143 = _ans_19_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_144 = _ans_19_leadingZeros_T_93[46] ? 6'h2e : _ans_19_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_145 = _ans_19_leadingZeros_T_93[45] ? 6'h2d : _ans_19_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_146 = _ans_19_leadingZeros_T_93[44] ? 6'h2c : _ans_19_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_147 = _ans_19_leadingZeros_T_93[43] ? 6'h2b : _ans_19_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_148 = _ans_19_leadingZeros_T_93[42] ? 6'h2a : _ans_19_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_149 = _ans_19_leadingZeros_T_93[41] ? 6'h29 : _ans_19_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_150 = _ans_19_leadingZeros_T_93[40] ? 6'h28 : _ans_19_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_151 = _ans_19_leadingZeros_T_93[39] ? 6'h27 : _ans_19_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_152 = _ans_19_leadingZeros_T_93[38] ? 6'h26 : _ans_19_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_153 = _ans_19_leadingZeros_T_93[37] ? 6'h25 : _ans_19_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_154 = _ans_19_leadingZeros_T_93[36] ? 6'h24 : _ans_19_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_155 = _ans_19_leadingZeros_T_93[35] ? 6'h23 : _ans_19_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_156 = _ans_19_leadingZeros_T_93[34] ? 6'h22 : _ans_19_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_157 = _ans_19_leadingZeros_T_93[33] ? 6'h21 : _ans_19_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_158 = _ans_19_leadingZeros_T_93[32] ? 6'h20 : _ans_19_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_159 = _ans_19_leadingZeros_T_93[31] ? 6'h1f : _ans_19_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_160 = _ans_19_leadingZeros_T_93[30] ? 6'h1e : _ans_19_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_161 = _ans_19_leadingZeros_T_93[29] ? 6'h1d : _ans_19_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_162 = _ans_19_leadingZeros_T_93[28] ? 6'h1c : _ans_19_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_163 = _ans_19_leadingZeros_T_93[27] ? 6'h1b : _ans_19_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_164 = _ans_19_leadingZeros_T_93[26] ? 6'h1a : _ans_19_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_165 = _ans_19_leadingZeros_T_93[25] ? 6'h19 : _ans_19_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_166 = _ans_19_leadingZeros_T_93[24] ? 6'h18 : _ans_19_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_167 = _ans_19_leadingZeros_T_93[23] ? 6'h17 : _ans_19_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_168 = _ans_19_leadingZeros_T_93[22] ? 6'h16 : _ans_19_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_169 = _ans_19_leadingZeros_T_93[21] ? 6'h15 : _ans_19_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_170 = _ans_19_leadingZeros_T_93[20] ? 6'h14 : _ans_19_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_171 = _ans_19_leadingZeros_T_93[19] ? 6'h13 : _ans_19_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_172 = _ans_19_leadingZeros_T_93[18] ? 6'h12 : _ans_19_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_173 = _ans_19_leadingZeros_T_93[17] ? 6'h11 : _ans_19_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_174 = _ans_19_leadingZeros_T_93[16] ? 6'h10 : _ans_19_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_175 = _ans_19_leadingZeros_T_93[15] ? 6'hf : _ans_19_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_176 = _ans_19_leadingZeros_T_93[14] ? 6'he : _ans_19_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_177 = _ans_19_leadingZeros_T_93[13] ? 6'hd : _ans_19_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_178 = _ans_19_leadingZeros_T_93[12] ? 6'hc : _ans_19_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_179 = _ans_19_leadingZeros_T_93[11] ? 6'hb : _ans_19_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_180 = _ans_19_leadingZeros_T_93[10] ? 6'ha : _ans_19_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_181 = _ans_19_leadingZeros_T_93[9] ? 6'h9 : _ans_19_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_182 = _ans_19_leadingZeros_T_93[8] ? 6'h8 : _ans_19_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_183 = _ans_19_leadingZeros_T_93[7] ? 6'h7 : _ans_19_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_184 = _ans_19_leadingZeros_T_93[6] ? 6'h6 : _ans_19_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_185 = _ans_19_leadingZeros_T_93[5] ? 6'h5 : _ans_19_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_186 = _ans_19_leadingZeros_T_93[4] ? 6'h4 : _ans_19_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_187 = _ans_19_leadingZeros_T_93[3] ? 6'h3 : _ans_19_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_188 = _ans_19_leadingZeros_T_93[2] ? 6'h2 : _ans_19_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_leadingZeros_T_189 = _ans_19_leadingZeros_T_93[1] ? 6'h1 : _ans_19_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_19_leadingZeros = _ans_19_leadingZeros_T_93[0] ? 6'h0 : _ans_19_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_19_expRaw_T_1 = 6'h1f - ans_19_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_19_expRaw = ans_19_isZero ? 6'h0 : _ans_19_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_19_shiftAmt_T_2 = ans_19_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_19_shiftAmt = ans_19_expRaw > 6'h3 ? _ans_19_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_19_mantissaRaw_T = ans_19_absClipped >> ans_19_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_19_mantissaRaw = _ans_19_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_19_mantissa = ans_19_expRaw >= 6'h3 ? ans_19_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_19_expAdjusted = ans_19_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_19_exp_T_4 = ans_19_expAdjusted > 7'hf ? 4'hf : ans_19_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_19_exp = ans_19_isZero ? 4'h0 : _ans_19_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_19_fp8 = {ans_19_clippedX[31],ans_19_exp,ans_19_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_20 = {24'h0,linear_bias_20}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_20 = tempSum_20 + biasExtended_20; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_20_sign = sum32_20[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_20_absX_T = ~sum32_20; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_20_absX_T_2 = _ans_20_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_20_absX = ans_20_sign ? _ans_20_absX_T_2 : sum32_20; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_20_shiftedX_T_1 = _GEN_14432 - ans_20_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_20_shiftedX_T_3 = ans_20_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_20_shiftedX = ans_20_sign ? _ans_20_shiftedX_T_1 : _ans_20_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_20_scaledX_T_1 = ans_20_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_20_scaledX = _ans_20_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_20_clippedX_T_2 = ans_20_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_20_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_20_clippedX = ans_20_scaledX > 49'h1c0 ? 49'h1c0 : _ans_20_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_20_absClipped_T_1 = ~ans_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_20_absClipped_T_3 = _ans_20_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_20_absClipped = ans_20_clippedX[31] ? _ans_20_absClipped_T_3 : ans_20_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_20_isZero = ans_20_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39934 = {{16'd0}, ans_20_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_4 = _GEN_39934 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_6 = {ans_20_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_8 = _ans_20_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_9 = _ans_20_leadingZeros_T_4 | _ans_20_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39935 = {{8'd0}, _ans_20_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_14 = _GEN_39935 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_16 = {_ans_20_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_18 = _ans_20_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_19 = _ans_20_leadingZeros_T_14 | _ans_20_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39936 = {{4'd0}, _ans_20_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_24 = _GEN_39936 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_26 = {_ans_20_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_28 = _ans_20_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_29 = _ans_20_leadingZeros_T_24 | _ans_20_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39937 = {{2'd0}, _ans_20_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_34 = _GEN_39937 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_36 = {_ans_20_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_38 = _ans_20_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_39 = _ans_20_leadingZeros_T_34 | _ans_20_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39938 = {{1'd0}, _ans_20_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_44 = _GEN_39938 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_46 = {_ans_20_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_48 = _ans_20_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_20_leadingZeros_T_49 = _ans_20_leadingZeros_T_44 | _ans_20_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39939 = {{8'd0}, ans_20_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_55 = _GEN_39939 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_57 = {ans_20_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_59 = _ans_20_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_60 = _ans_20_leadingZeros_T_55 | _ans_20_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39940 = {{4'd0}, _ans_20_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_65 = _GEN_39940 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_67 = {_ans_20_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_69 = _ans_20_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_70 = _ans_20_leadingZeros_T_65 | _ans_20_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39941 = {{2'd0}, _ans_20_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_75 = _GEN_39941 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_77 = {_ans_20_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_79 = _ans_20_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_80 = _ans_20_leadingZeros_T_75 | _ans_20_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39942 = {{1'd0}, _ans_20_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_85 = _GEN_39942 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_87 = {_ans_20_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_89 = _ans_20_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_20_leadingZeros_T_90 = _ans_20_leadingZeros_T_85 | _ans_20_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_20_leadingZeros_T_93 = {_ans_20_leadingZeros_T_49,_ans_20_leadingZeros_T_90,ans_20_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_20_leadingZeros_T_143 = _ans_20_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_144 = _ans_20_leadingZeros_T_93[46] ? 6'h2e : _ans_20_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_145 = _ans_20_leadingZeros_T_93[45] ? 6'h2d : _ans_20_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_146 = _ans_20_leadingZeros_T_93[44] ? 6'h2c : _ans_20_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_147 = _ans_20_leadingZeros_T_93[43] ? 6'h2b : _ans_20_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_148 = _ans_20_leadingZeros_T_93[42] ? 6'h2a : _ans_20_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_149 = _ans_20_leadingZeros_T_93[41] ? 6'h29 : _ans_20_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_150 = _ans_20_leadingZeros_T_93[40] ? 6'h28 : _ans_20_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_151 = _ans_20_leadingZeros_T_93[39] ? 6'h27 : _ans_20_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_152 = _ans_20_leadingZeros_T_93[38] ? 6'h26 : _ans_20_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_153 = _ans_20_leadingZeros_T_93[37] ? 6'h25 : _ans_20_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_154 = _ans_20_leadingZeros_T_93[36] ? 6'h24 : _ans_20_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_155 = _ans_20_leadingZeros_T_93[35] ? 6'h23 : _ans_20_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_156 = _ans_20_leadingZeros_T_93[34] ? 6'h22 : _ans_20_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_157 = _ans_20_leadingZeros_T_93[33] ? 6'h21 : _ans_20_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_158 = _ans_20_leadingZeros_T_93[32] ? 6'h20 : _ans_20_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_159 = _ans_20_leadingZeros_T_93[31] ? 6'h1f : _ans_20_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_160 = _ans_20_leadingZeros_T_93[30] ? 6'h1e : _ans_20_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_161 = _ans_20_leadingZeros_T_93[29] ? 6'h1d : _ans_20_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_162 = _ans_20_leadingZeros_T_93[28] ? 6'h1c : _ans_20_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_163 = _ans_20_leadingZeros_T_93[27] ? 6'h1b : _ans_20_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_164 = _ans_20_leadingZeros_T_93[26] ? 6'h1a : _ans_20_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_165 = _ans_20_leadingZeros_T_93[25] ? 6'h19 : _ans_20_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_166 = _ans_20_leadingZeros_T_93[24] ? 6'h18 : _ans_20_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_167 = _ans_20_leadingZeros_T_93[23] ? 6'h17 : _ans_20_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_168 = _ans_20_leadingZeros_T_93[22] ? 6'h16 : _ans_20_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_169 = _ans_20_leadingZeros_T_93[21] ? 6'h15 : _ans_20_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_170 = _ans_20_leadingZeros_T_93[20] ? 6'h14 : _ans_20_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_171 = _ans_20_leadingZeros_T_93[19] ? 6'h13 : _ans_20_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_172 = _ans_20_leadingZeros_T_93[18] ? 6'h12 : _ans_20_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_173 = _ans_20_leadingZeros_T_93[17] ? 6'h11 : _ans_20_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_174 = _ans_20_leadingZeros_T_93[16] ? 6'h10 : _ans_20_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_175 = _ans_20_leadingZeros_T_93[15] ? 6'hf : _ans_20_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_176 = _ans_20_leadingZeros_T_93[14] ? 6'he : _ans_20_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_177 = _ans_20_leadingZeros_T_93[13] ? 6'hd : _ans_20_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_178 = _ans_20_leadingZeros_T_93[12] ? 6'hc : _ans_20_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_179 = _ans_20_leadingZeros_T_93[11] ? 6'hb : _ans_20_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_180 = _ans_20_leadingZeros_T_93[10] ? 6'ha : _ans_20_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_181 = _ans_20_leadingZeros_T_93[9] ? 6'h9 : _ans_20_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_182 = _ans_20_leadingZeros_T_93[8] ? 6'h8 : _ans_20_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_183 = _ans_20_leadingZeros_T_93[7] ? 6'h7 : _ans_20_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_184 = _ans_20_leadingZeros_T_93[6] ? 6'h6 : _ans_20_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_185 = _ans_20_leadingZeros_T_93[5] ? 6'h5 : _ans_20_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_186 = _ans_20_leadingZeros_T_93[4] ? 6'h4 : _ans_20_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_187 = _ans_20_leadingZeros_T_93[3] ? 6'h3 : _ans_20_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_188 = _ans_20_leadingZeros_T_93[2] ? 6'h2 : _ans_20_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_leadingZeros_T_189 = _ans_20_leadingZeros_T_93[1] ? 6'h1 : _ans_20_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_20_leadingZeros = _ans_20_leadingZeros_T_93[0] ? 6'h0 : _ans_20_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_20_expRaw_T_1 = 6'h1f - ans_20_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_20_expRaw = ans_20_isZero ? 6'h0 : _ans_20_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_20_shiftAmt_T_2 = ans_20_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_20_shiftAmt = ans_20_expRaw > 6'h3 ? _ans_20_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_20_mantissaRaw_T = ans_20_absClipped >> ans_20_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_20_mantissaRaw = _ans_20_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_20_mantissa = ans_20_expRaw >= 6'h3 ? ans_20_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_20_expAdjusted = ans_20_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_20_exp_T_4 = ans_20_expAdjusted > 7'hf ? 4'hf : ans_20_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_20_exp = ans_20_isZero ? 4'h0 : _ans_20_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_20_fp8 = {ans_20_clippedX[31],ans_20_exp,ans_20_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_21 = {24'h0,linear_bias_21}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_21 = tempSum_21 + biasExtended_21; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_21_sign = sum32_21[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_21_absX_T = ~sum32_21; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_21_absX_T_2 = _ans_21_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_21_absX = ans_21_sign ? _ans_21_absX_T_2 : sum32_21; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_21_shiftedX_T_1 = _GEN_14432 - ans_21_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_21_shiftedX_T_3 = ans_21_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_21_shiftedX = ans_21_sign ? _ans_21_shiftedX_T_1 : _ans_21_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_21_scaledX_T_1 = ans_21_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_21_scaledX = _ans_21_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_21_clippedX_T_2 = ans_21_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_21_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_21_clippedX = ans_21_scaledX > 49'h1c0 ? 49'h1c0 : _ans_21_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_21_absClipped_T_1 = ~ans_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_21_absClipped_T_3 = _ans_21_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_21_absClipped = ans_21_clippedX[31] ? _ans_21_absClipped_T_3 : ans_21_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_21_isZero = ans_21_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39945 = {{16'd0}, ans_21_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_4 = _GEN_39945 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_6 = {ans_21_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_8 = _ans_21_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_9 = _ans_21_leadingZeros_T_4 | _ans_21_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39946 = {{8'd0}, _ans_21_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_14 = _GEN_39946 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_16 = {_ans_21_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_18 = _ans_21_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_19 = _ans_21_leadingZeros_T_14 | _ans_21_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39947 = {{4'd0}, _ans_21_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_24 = _GEN_39947 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_26 = {_ans_21_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_28 = _ans_21_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_29 = _ans_21_leadingZeros_T_24 | _ans_21_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39948 = {{2'd0}, _ans_21_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_34 = _GEN_39948 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_36 = {_ans_21_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_38 = _ans_21_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_39 = _ans_21_leadingZeros_T_34 | _ans_21_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39949 = {{1'd0}, _ans_21_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_44 = _GEN_39949 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_46 = {_ans_21_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_48 = _ans_21_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_21_leadingZeros_T_49 = _ans_21_leadingZeros_T_44 | _ans_21_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39950 = {{8'd0}, ans_21_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_55 = _GEN_39950 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_57 = {ans_21_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_59 = _ans_21_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_60 = _ans_21_leadingZeros_T_55 | _ans_21_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39951 = {{4'd0}, _ans_21_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_65 = _GEN_39951 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_67 = {_ans_21_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_69 = _ans_21_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_70 = _ans_21_leadingZeros_T_65 | _ans_21_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39952 = {{2'd0}, _ans_21_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_75 = _GEN_39952 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_77 = {_ans_21_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_79 = _ans_21_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_80 = _ans_21_leadingZeros_T_75 | _ans_21_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39953 = {{1'd0}, _ans_21_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_85 = _GEN_39953 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_87 = {_ans_21_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_89 = _ans_21_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_21_leadingZeros_T_90 = _ans_21_leadingZeros_T_85 | _ans_21_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_21_leadingZeros_T_93 = {_ans_21_leadingZeros_T_49,_ans_21_leadingZeros_T_90,ans_21_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_21_leadingZeros_T_143 = _ans_21_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_144 = _ans_21_leadingZeros_T_93[46] ? 6'h2e : _ans_21_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_145 = _ans_21_leadingZeros_T_93[45] ? 6'h2d : _ans_21_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_146 = _ans_21_leadingZeros_T_93[44] ? 6'h2c : _ans_21_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_147 = _ans_21_leadingZeros_T_93[43] ? 6'h2b : _ans_21_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_148 = _ans_21_leadingZeros_T_93[42] ? 6'h2a : _ans_21_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_149 = _ans_21_leadingZeros_T_93[41] ? 6'h29 : _ans_21_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_150 = _ans_21_leadingZeros_T_93[40] ? 6'h28 : _ans_21_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_151 = _ans_21_leadingZeros_T_93[39] ? 6'h27 : _ans_21_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_152 = _ans_21_leadingZeros_T_93[38] ? 6'h26 : _ans_21_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_153 = _ans_21_leadingZeros_T_93[37] ? 6'h25 : _ans_21_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_154 = _ans_21_leadingZeros_T_93[36] ? 6'h24 : _ans_21_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_155 = _ans_21_leadingZeros_T_93[35] ? 6'h23 : _ans_21_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_156 = _ans_21_leadingZeros_T_93[34] ? 6'h22 : _ans_21_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_157 = _ans_21_leadingZeros_T_93[33] ? 6'h21 : _ans_21_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_158 = _ans_21_leadingZeros_T_93[32] ? 6'h20 : _ans_21_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_159 = _ans_21_leadingZeros_T_93[31] ? 6'h1f : _ans_21_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_160 = _ans_21_leadingZeros_T_93[30] ? 6'h1e : _ans_21_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_161 = _ans_21_leadingZeros_T_93[29] ? 6'h1d : _ans_21_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_162 = _ans_21_leadingZeros_T_93[28] ? 6'h1c : _ans_21_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_163 = _ans_21_leadingZeros_T_93[27] ? 6'h1b : _ans_21_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_164 = _ans_21_leadingZeros_T_93[26] ? 6'h1a : _ans_21_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_165 = _ans_21_leadingZeros_T_93[25] ? 6'h19 : _ans_21_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_166 = _ans_21_leadingZeros_T_93[24] ? 6'h18 : _ans_21_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_167 = _ans_21_leadingZeros_T_93[23] ? 6'h17 : _ans_21_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_168 = _ans_21_leadingZeros_T_93[22] ? 6'h16 : _ans_21_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_169 = _ans_21_leadingZeros_T_93[21] ? 6'h15 : _ans_21_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_170 = _ans_21_leadingZeros_T_93[20] ? 6'h14 : _ans_21_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_171 = _ans_21_leadingZeros_T_93[19] ? 6'h13 : _ans_21_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_172 = _ans_21_leadingZeros_T_93[18] ? 6'h12 : _ans_21_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_173 = _ans_21_leadingZeros_T_93[17] ? 6'h11 : _ans_21_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_174 = _ans_21_leadingZeros_T_93[16] ? 6'h10 : _ans_21_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_175 = _ans_21_leadingZeros_T_93[15] ? 6'hf : _ans_21_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_176 = _ans_21_leadingZeros_T_93[14] ? 6'he : _ans_21_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_177 = _ans_21_leadingZeros_T_93[13] ? 6'hd : _ans_21_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_178 = _ans_21_leadingZeros_T_93[12] ? 6'hc : _ans_21_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_179 = _ans_21_leadingZeros_T_93[11] ? 6'hb : _ans_21_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_180 = _ans_21_leadingZeros_T_93[10] ? 6'ha : _ans_21_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_181 = _ans_21_leadingZeros_T_93[9] ? 6'h9 : _ans_21_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_182 = _ans_21_leadingZeros_T_93[8] ? 6'h8 : _ans_21_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_183 = _ans_21_leadingZeros_T_93[7] ? 6'h7 : _ans_21_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_184 = _ans_21_leadingZeros_T_93[6] ? 6'h6 : _ans_21_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_185 = _ans_21_leadingZeros_T_93[5] ? 6'h5 : _ans_21_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_186 = _ans_21_leadingZeros_T_93[4] ? 6'h4 : _ans_21_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_187 = _ans_21_leadingZeros_T_93[3] ? 6'h3 : _ans_21_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_188 = _ans_21_leadingZeros_T_93[2] ? 6'h2 : _ans_21_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_leadingZeros_T_189 = _ans_21_leadingZeros_T_93[1] ? 6'h1 : _ans_21_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_21_leadingZeros = _ans_21_leadingZeros_T_93[0] ? 6'h0 : _ans_21_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_21_expRaw_T_1 = 6'h1f - ans_21_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_21_expRaw = ans_21_isZero ? 6'h0 : _ans_21_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_21_shiftAmt_T_2 = ans_21_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_21_shiftAmt = ans_21_expRaw > 6'h3 ? _ans_21_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_21_mantissaRaw_T = ans_21_absClipped >> ans_21_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_21_mantissaRaw = _ans_21_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_21_mantissa = ans_21_expRaw >= 6'h3 ? ans_21_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_21_expAdjusted = ans_21_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_21_exp_T_4 = ans_21_expAdjusted > 7'hf ? 4'hf : ans_21_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_21_exp = ans_21_isZero ? 4'h0 : _ans_21_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_21_fp8 = {ans_21_clippedX[31],ans_21_exp,ans_21_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_22 = {24'h0,linear_bias_22}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_22 = tempSum_22 + biasExtended_22; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_22_sign = sum32_22[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_22_absX_T = ~sum32_22; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_22_absX_T_2 = _ans_22_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_22_absX = ans_22_sign ? _ans_22_absX_T_2 : sum32_22; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_22_shiftedX_T_1 = _GEN_14432 - ans_22_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_22_shiftedX_T_3 = ans_22_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_22_shiftedX = ans_22_sign ? _ans_22_shiftedX_T_1 : _ans_22_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_22_scaledX_T_1 = ans_22_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_22_scaledX = _ans_22_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_22_clippedX_T_2 = ans_22_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_22_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_22_clippedX = ans_22_scaledX > 49'h1c0 ? 49'h1c0 : _ans_22_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_22_absClipped_T_1 = ~ans_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_22_absClipped_T_3 = _ans_22_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_22_absClipped = ans_22_clippedX[31] ? _ans_22_absClipped_T_3 : ans_22_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_22_isZero = ans_22_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39956 = {{16'd0}, ans_22_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_4 = _GEN_39956 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_6 = {ans_22_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_8 = _ans_22_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_9 = _ans_22_leadingZeros_T_4 | _ans_22_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39957 = {{8'd0}, _ans_22_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_14 = _GEN_39957 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_16 = {_ans_22_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_18 = _ans_22_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_19 = _ans_22_leadingZeros_T_14 | _ans_22_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39958 = {{4'd0}, _ans_22_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_24 = _GEN_39958 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_26 = {_ans_22_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_28 = _ans_22_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_29 = _ans_22_leadingZeros_T_24 | _ans_22_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39959 = {{2'd0}, _ans_22_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_34 = _GEN_39959 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_36 = {_ans_22_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_38 = _ans_22_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_39 = _ans_22_leadingZeros_T_34 | _ans_22_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39960 = {{1'd0}, _ans_22_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_44 = _GEN_39960 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_46 = {_ans_22_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_48 = _ans_22_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_22_leadingZeros_T_49 = _ans_22_leadingZeros_T_44 | _ans_22_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39961 = {{8'd0}, ans_22_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_55 = _GEN_39961 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_57 = {ans_22_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_59 = _ans_22_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_60 = _ans_22_leadingZeros_T_55 | _ans_22_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39962 = {{4'd0}, _ans_22_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_65 = _GEN_39962 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_67 = {_ans_22_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_69 = _ans_22_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_70 = _ans_22_leadingZeros_T_65 | _ans_22_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39963 = {{2'd0}, _ans_22_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_75 = _GEN_39963 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_77 = {_ans_22_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_79 = _ans_22_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_80 = _ans_22_leadingZeros_T_75 | _ans_22_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39964 = {{1'd0}, _ans_22_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_85 = _GEN_39964 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_87 = {_ans_22_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_89 = _ans_22_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_22_leadingZeros_T_90 = _ans_22_leadingZeros_T_85 | _ans_22_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_22_leadingZeros_T_93 = {_ans_22_leadingZeros_T_49,_ans_22_leadingZeros_T_90,ans_22_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_22_leadingZeros_T_143 = _ans_22_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_144 = _ans_22_leadingZeros_T_93[46] ? 6'h2e : _ans_22_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_145 = _ans_22_leadingZeros_T_93[45] ? 6'h2d : _ans_22_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_146 = _ans_22_leadingZeros_T_93[44] ? 6'h2c : _ans_22_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_147 = _ans_22_leadingZeros_T_93[43] ? 6'h2b : _ans_22_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_148 = _ans_22_leadingZeros_T_93[42] ? 6'h2a : _ans_22_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_149 = _ans_22_leadingZeros_T_93[41] ? 6'h29 : _ans_22_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_150 = _ans_22_leadingZeros_T_93[40] ? 6'h28 : _ans_22_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_151 = _ans_22_leadingZeros_T_93[39] ? 6'h27 : _ans_22_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_152 = _ans_22_leadingZeros_T_93[38] ? 6'h26 : _ans_22_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_153 = _ans_22_leadingZeros_T_93[37] ? 6'h25 : _ans_22_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_154 = _ans_22_leadingZeros_T_93[36] ? 6'h24 : _ans_22_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_155 = _ans_22_leadingZeros_T_93[35] ? 6'h23 : _ans_22_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_156 = _ans_22_leadingZeros_T_93[34] ? 6'h22 : _ans_22_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_157 = _ans_22_leadingZeros_T_93[33] ? 6'h21 : _ans_22_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_158 = _ans_22_leadingZeros_T_93[32] ? 6'h20 : _ans_22_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_159 = _ans_22_leadingZeros_T_93[31] ? 6'h1f : _ans_22_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_160 = _ans_22_leadingZeros_T_93[30] ? 6'h1e : _ans_22_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_161 = _ans_22_leadingZeros_T_93[29] ? 6'h1d : _ans_22_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_162 = _ans_22_leadingZeros_T_93[28] ? 6'h1c : _ans_22_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_163 = _ans_22_leadingZeros_T_93[27] ? 6'h1b : _ans_22_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_164 = _ans_22_leadingZeros_T_93[26] ? 6'h1a : _ans_22_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_165 = _ans_22_leadingZeros_T_93[25] ? 6'h19 : _ans_22_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_166 = _ans_22_leadingZeros_T_93[24] ? 6'h18 : _ans_22_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_167 = _ans_22_leadingZeros_T_93[23] ? 6'h17 : _ans_22_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_168 = _ans_22_leadingZeros_T_93[22] ? 6'h16 : _ans_22_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_169 = _ans_22_leadingZeros_T_93[21] ? 6'h15 : _ans_22_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_170 = _ans_22_leadingZeros_T_93[20] ? 6'h14 : _ans_22_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_171 = _ans_22_leadingZeros_T_93[19] ? 6'h13 : _ans_22_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_172 = _ans_22_leadingZeros_T_93[18] ? 6'h12 : _ans_22_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_173 = _ans_22_leadingZeros_T_93[17] ? 6'h11 : _ans_22_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_174 = _ans_22_leadingZeros_T_93[16] ? 6'h10 : _ans_22_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_175 = _ans_22_leadingZeros_T_93[15] ? 6'hf : _ans_22_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_176 = _ans_22_leadingZeros_T_93[14] ? 6'he : _ans_22_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_177 = _ans_22_leadingZeros_T_93[13] ? 6'hd : _ans_22_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_178 = _ans_22_leadingZeros_T_93[12] ? 6'hc : _ans_22_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_179 = _ans_22_leadingZeros_T_93[11] ? 6'hb : _ans_22_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_180 = _ans_22_leadingZeros_T_93[10] ? 6'ha : _ans_22_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_181 = _ans_22_leadingZeros_T_93[9] ? 6'h9 : _ans_22_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_182 = _ans_22_leadingZeros_T_93[8] ? 6'h8 : _ans_22_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_183 = _ans_22_leadingZeros_T_93[7] ? 6'h7 : _ans_22_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_184 = _ans_22_leadingZeros_T_93[6] ? 6'h6 : _ans_22_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_185 = _ans_22_leadingZeros_T_93[5] ? 6'h5 : _ans_22_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_186 = _ans_22_leadingZeros_T_93[4] ? 6'h4 : _ans_22_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_187 = _ans_22_leadingZeros_T_93[3] ? 6'h3 : _ans_22_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_188 = _ans_22_leadingZeros_T_93[2] ? 6'h2 : _ans_22_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_leadingZeros_T_189 = _ans_22_leadingZeros_T_93[1] ? 6'h1 : _ans_22_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_22_leadingZeros = _ans_22_leadingZeros_T_93[0] ? 6'h0 : _ans_22_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_22_expRaw_T_1 = 6'h1f - ans_22_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_22_expRaw = ans_22_isZero ? 6'h0 : _ans_22_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_22_shiftAmt_T_2 = ans_22_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_22_shiftAmt = ans_22_expRaw > 6'h3 ? _ans_22_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_22_mantissaRaw_T = ans_22_absClipped >> ans_22_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_22_mantissaRaw = _ans_22_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_22_mantissa = ans_22_expRaw >= 6'h3 ? ans_22_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_22_expAdjusted = ans_22_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_22_exp_T_4 = ans_22_expAdjusted > 7'hf ? 4'hf : ans_22_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_22_exp = ans_22_isZero ? 4'h0 : _ans_22_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_22_fp8 = {ans_22_clippedX[31],ans_22_exp,ans_22_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_23 = {24'h0,linear_bias_23}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_23 = tempSum_23 + biasExtended_23; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_23_sign = sum32_23[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_23_absX_T = ~sum32_23; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_23_absX_T_2 = _ans_23_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_23_absX = ans_23_sign ? _ans_23_absX_T_2 : sum32_23; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_23_shiftedX_T_1 = _GEN_14432 - ans_23_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_23_shiftedX_T_3 = ans_23_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_23_shiftedX = ans_23_sign ? _ans_23_shiftedX_T_1 : _ans_23_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_23_scaledX_T_1 = ans_23_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_23_scaledX = _ans_23_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_23_clippedX_T_2 = ans_23_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_23_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_23_clippedX = ans_23_scaledX > 49'h1c0 ? 49'h1c0 : _ans_23_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_23_absClipped_T_1 = ~ans_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_23_absClipped_T_3 = _ans_23_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_23_absClipped = ans_23_clippedX[31] ? _ans_23_absClipped_T_3 : ans_23_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_23_isZero = ans_23_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39967 = {{16'd0}, ans_23_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_4 = _GEN_39967 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_6 = {ans_23_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_8 = _ans_23_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_9 = _ans_23_leadingZeros_T_4 | _ans_23_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39968 = {{8'd0}, _ans_23_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_14 = _GEN_39968 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_16 = {_ans_23_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_18 = _ans_23_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_19 = _ans_23_leadingZeros_T_14 | _ans_23_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39969 = {{4'd0}, _ans_23_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_24 = _GEN_39969 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_26 = {_ans_23_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_28 = _ans_23_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_29 = _ans_23_leadingZeros_T_24 | _ans_23_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39970 = {{2'd0}, _ans_23_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_34 = _GEN_39970 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_36 = {_ans_23_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_38 = _ans_23_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_39 = _ans_23_leadingZeros_T_34 | _ans_23_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39971 = {{1'd0}, _ans_23_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_44 = _GEN_39971 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_46 = {_ans_23_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_48 = _ans_23_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_23_leadingZeros_T_49 = _ans_23_leadingZeros_T_44 | _ans_23_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39972 = {{8'd0}, ans_23_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_55 = _GEN_39972 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_57 = {ans_23_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_59 = _ans_23_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_60 = _ans_23_leadingZeros_T_55 | _ans_23_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39973 = {{4'd0}, _ans_23_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_65 = _GEN_39973 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_67 = {_ans_23_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_69 = _ans_23_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_70 = _ans_23_leadingZeros_T_65 | _ans_23_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39974 = {{2'd0}, _ans_23_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_75 = _GEN_39974 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_77 = {_ans_23_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_79 = _ans_23_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_80 = _ans_23_leadingZeros_T_75 | _ans_23_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39975 = {{1'd0}, _ans_23_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_85 = _GEN_39975 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_87 = {_ans_23_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_89 = _ans_23_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_23_leadingZeros_T_90 = _ans_23_leadingZeros_T_85 | _ans_23_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_23_leadingZeros_T_93 = {_ans_23_leadingZeros_T_49,_ans_23_leadingZeros_T_90,ans_23_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_23_leadingZeros_T_143 = _ans_23_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_144 = _ans_23_leadingZeros_T_93[46] ? 6'h2e : _ans_23_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_145 = _ans_23_leadingZeros_T_93[45] ? 6'h2d : _ans_23_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_146 = _ans_23_leadingZeros_T_93[44] ? 6'h2c : _ans_23_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_147 = _ans_23_leadingZeros_T_93[43] ? 6'h2b : _ans_23_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_148 = _ans_23_leadingZeros_T_93[42] ? 6'h2a : _ans_23_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_149 = _ans_23_leadingZeros_T_93[41] ? 6'h29 : _ans_23_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_150 = _ans_23_leadingZeros_T_93[40] ? 6'h28 : _ans_23_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_151 = _ans_23_leadingZeros_T_93[39] ? 6'h27 : _ans_23_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_152 = _ans_23_leadingZeros_T_93[38] ? 6'h26 : _ans_23_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_153 = _ans_23_leadingZeros_T_93[37] ? 6'h25 : _ans_23_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_154 = _ans_23_leadingZeros_T_93[36] ? 6'h24 : _ans_23_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_155 = _ans_23_leadingZeros_T_93[35] ? 6'h23 : _ans_23_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_156 = _ans_23_leadingZeros_T_93[34] ? 6'h22 : _ans_23_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_157 = _ans_23_leadingZeros_T_93[33] ? 6'h21 : _ans_23_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_158 = _ans_23_leadingZeros_T_93[32] ? 6'h20 : _ans_23_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_159 = _ans_23_leadingZeros_T_93[31] ? 6'h1f : _ans_23_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_160 = _ans_23_leadingZeros_T_93[30] ? 6'h1e : _ans_23_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_161 = _ans_23_leadingZeros_T_93[29] ? 6'h1d : _ans_23_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_162 = _ans_23_leadingZeros_T_93[28] ? 6'h1c : _ans_23_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_163 = _ans_23_leadingZeros_T_93[27] ? 6'h1b : _ans_23_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_164 = _ans_23_leadingZeros_T_93[26] ? 6'h1a : _ans_23_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_165 = _ans_23_leadingZeros_T_93[25] ? 6'h19 : _ans_23_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_166 = _ans_23_leadingZeros_T_93[24] ? 6'h18 : _ans_23_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_167 = _ans_23_leadingZeros_T_93[23] ? 6'h17 : _ans_23_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_168 = _ans_23_leadingZeros_T_93[22] ? 6'h16 : _ans_23_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_169 = _ans_23_leadingZeros_T_93[21] ? 6'h15 : _ans_23_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_170 = _ans_23_leadingZeros_T_93[20] ? 6'h14 : _ans_23_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_171 = _ans_23_leadingZeros_T_93[19] ? 6'h13 : _ans_23_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_172 = _ans_23_leadingZeros_T_93[18] ? 6'h12 : _ans_23_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_173 = _ans_23_leadingZeros_T_93[17] ? 6'h11 : _ans_23_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_174 = _ans_23_leadingZeros_T_93[16] ? 6'h10 : _ans_23_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_175 = _ans_23_leadingZeros_T_93[15] ? 6'hf : _ans_23_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_176 = _ans_23_leadingZeros_T_93[14] ? 6'he : _ans_23_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_177 = _ans_23_leadingZeros_T_93[13] ? 6'hd : _ans_23_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_178 = _ans_23_leadingZeros_T_93[12] ? 6'hc : _ans_23_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_179 = _ans_23_leadingZeros_T_93[11] ? 6'hb : _ans_23_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_180 = _ans_23_leadingZeros_T_93[10] ? 6'ha : _ans_23_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_181 = _ans_23_leadingZeros_T_93[9] ? 6'h9 : _ans_23_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_182 = _ans_23_leadingZeros_T_93[8] ? 6'h8 : _ans_23_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_183 = _ans_23_leadingZeros_T_93[7] ? 6'h7 : _ans_23_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_184 = _ans_23_leadingZeros_T_93[6] ? 6'h6 : _ans_23_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_185 = _ans_23_leadingZeros_T_93[5] ? 6'h5 : _ans_23_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_186 = _ans_23_leadingZeros_T_93[4] ? 6'h4 : _ans_23_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_187 = _ans_23_leadingZeros_T_93[3] ? 6'h3 : _ans_23_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_188 = _ans_23_leadingZeros_T_93[2] ? 6'h2 : _ans_23_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_leadingZeros_T_189 = _ans_23_leadingZeros_T_93[1] ? 6'h1 : _ans_23_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_23_leadingZeros = _ans_23_leadingZeros_T_93[0] ? 6'h0 : _ans_23_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_23_expRaw_T_1 = 6'h1f - ans_23_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_23_expRaw = ans_23_isZero ? 6'h0 : _ans_23_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_23_shiftAmt_T_2 = ans_23_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_23_shiftAmt = ans_23_expRaw > 6'h3 ? _ans_23_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_23_mantissaRaw_T = ans_23_absClipped >> ans_23_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_23_mantissaRaw = _ans_23_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_23_mantissa = ans_23_expRaw >= 6'h3 ? ans_23_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_23_expAdjusted = ans_23_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_23_exp_T_4 = ans_23_expAdjusted > 7'hf ? 4'hf : ans_23_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_23_exp = ans_23_isZero ? 4'h0 : _ans_23_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_23_fp8 = {ans_23_clippedX[31],ans_23_exp,ans_23_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_24 = {24'h0,linear_bias_24}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_24 = tempSum_24 + biasExtended_24; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_24_sign = sum32_24[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_24_absX_T = ~sum32_24; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_24_absX_T_2 = _ans_24_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_24_absX = ans_24_sign ? _ans_24_absX_T_2 : sum32_24; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_24_shiftedX_T_1 = _GEN_14432 - ans_24_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_24_shiftedX_T_3 = ans_24_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_24_shiftedX = ans_24_sign ? _ans_24_shiftedX_T_1 : _ans_24_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_24_scaledX_T_1 = ans_24_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_24_scaledX = _ans_24_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_24_clippedX_T_2 = ans_24_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_24_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_24_clippedX = ans_24_scaledX > 49'h1c0 ? 49'h1c0 : _ans_24_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_24_absClipped_T_1 = ~ans_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_24_absClipped_T_3 = _ans_24_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_24_absClipped = ans_24_clippedX[31] ? _ans_24_absClipped_T_3 : ans_24_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_24_isZero = ans_24_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39978 = {{16'd0}, ans_24_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_4 = _GEN_39978 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_6 = {ans_24_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_8 = _ans_24_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_9 = _ans_24_leadingZeros_T_4 | _ans_24_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39979 = {{8'd0}, _ans_24_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_14 = _GEN_39979 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_16 = {_ans_24_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_18 = _ans_24_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_19 = _ans_24_leadingZeros_T_14 | _ans_24_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39980 = {{4'd0}, _ans_24_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_24 = _GEN_39980 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_26 = {_ans_24_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_28 = _ans_24_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_29 = _ans_24_leadingZeros_T_24 | _ans_24_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39981 = {{2'd0}, _ans_24_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_34 = _GEN_39981 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_36 = {_ans_24_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_38 = _ans_24_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_39 = _ans_24_leadingZeros_T_34 | _ans_24_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39982 = {{1'd0}, _ans_24_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_44 = _GEN_39982 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_46 = {_ans_24_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_48 = _ans_24_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_24_leadingZeros_T_49 = _ans_24_leadingZeros_T_44 | _ans_24_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39983 = {{8'd0}, ans_24_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_55 = _GEN_39983 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_57 = {ans_24_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_59 = _ans_24_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_60 = _ans_24_leadingZeros_T_55 | _ans_24_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39984 = {{4'd0}, _ans_24_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_65 = _GEN_39984 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_67 = {_ans_24_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_69 = _ans_24_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_70 = _ans_24_leadingZeros_T_65 | _ans_24_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39985 = {{2'd0}, _ans_24_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_75 = _GEN_39985 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_77 = {_ans_24_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_79 = _ans_24_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_80 = _ans_24_leadingZeros_T_75 | _ans_24_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39986 = {{1'd0}, _ans_24_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_85 = _GEN_39986 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_87 = {_ans_24_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_89 = _ans_24_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_24_leadingZeros_T_90 = _ans_24_leadingZeros_T_85 | _ans_24_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_24_leadingZeros_T_93 = {_ans_24_leadingZeros_T_49,_ans_24_leadingZeros_T_90,ans_24_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_24_leadingZeros_T_143 = _ans_24_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_144 = _ans_24_leadingZeros_T_93[46] ? 6'h2e : _ans_24_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_145 = _ans_24_leadingZeros_T_93[45] ? 6'h2d : _ans_24_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_146 = _ans_24_leadingZeros_T_93[44] ? 6'h2c : _ans_24_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_147 = _ans_24_leadingZeros_T_93[43] ? 6'h2b : _ans_24_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_148 = _ans_24_leadingZeros_T_93[42] ? 6'h2a : _ans_24_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_149 = _ans_24_leadingZeros_T_93[41] ? 6'h29 : _ans_24_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_150 = _ans_24_leadingZeros_T_93[40] ? 6'h28 : _ans_24_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_151 = _ans_24_leadingZeros_T_93[39] ? 6'h27 : _ans_24_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_152 = _ans_24_leadingZeros_T_93[38] ? 6'h26 : _ans_24_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_153 = _ans_24_leadingZeros_T_93[37] ? 6'h25 : _ans_24_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_154 = _ans_24_leadingZeros_T_93[36] ? 6'h24 : _ans_24_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_155 = _ans_24_leadingZeros_T_93[35] ? 6'h23 : _ans_24_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_156 = _ans_24_leadingZeros_T_93[34] ? 6'h22 : _ans_24_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_157 = _ans_24_leadingZeros_T_93[33] ? 6'h21 : _ans_24_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_158 = _ans_24_leadingZeros_T_93[32] ? 6'h20 : _ans_24_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_159 = _ans_24_leadingZeros_T_93[31] ? 6'h1f : _ans_24_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_160 = _ans_24_leadingZeros_T_93[30] ? 6'h1e : _ans_24_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_161 = _ans_24_leadingZeros_T_93[29] ? 6'h1d : _ans_24_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_162 = _ans_24_leadingZeros_T_93[28] ? 6'h1c : _ans_24_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_163 = _ans_24_leadingZeros_T_93[27] ? 6'h1b : _ans_24_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_164 = _ans_24_leadingZeros_T_93[26] ? 6'h1a : _ans_24_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_165 = _ans_24_leadingZeros_T_93[25] ? 6'h19 : _ans_24_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_166 = _ans_24_leadingZeros_T_93[24] ? 6'h18 : _ans_24_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_167 = _ans_24_leadingZeros_T_93[23] ? 6'h17 : _ans_24_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_168 = _ans_24_leadingZeros_T_93[22] ? 6'h16 : _ans_24_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_169 = _ans_24_leadingZeros_T_93[21] ? 6'h15 : _ans_24_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_170 = _ans_24_leadingZeros_T_93[20] ? 6'h14 : _ans_24_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_171 = _ans_24_leadingZeros_T_93[19] ? 6'h13 : _ans_24_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_172 = _ans_24_leadingZeros_T_93[18] ? 6'h12 : _ans_24_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_173 = _ans_24_leadingZeros_T_93[17] ? 6'h11 : _ans_24_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_174 = _ans_24_leadingZeros_T_93[16] ? 6'h10 : _ans_24_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_175 = _ans_24_leadingZeros_T_93[15] ? 6'hf : _ans_24_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_176 = _ans_24_leadingZeros_T_93[14] ? 6'he : _ans_24_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_177 = _ans_24_leadingZeros_T_93[13] ? 6'hd : _ans_24_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_178 = _ans_24_leadingZeros_T_93[12] ? 6'hc : _ans_24_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_179 = _ans_24_leadingZeros_T_93[11] ? 6'hb : _ans_24_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_180 = _ans_24_leadingZeros_T_93[10] ? 6'ha : _ans_24_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_181 = _ans_24_leadingZeros_T_93[9] ? 6'h9 : _ans_24_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_182 = _ans_24_leadingZeros_T_93[8] ? 6'h8 : _ans_24_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_183 = _ans_24_leadingZeros_T_93[7] ? 6'h7 : _ans_24_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_184 = _ans_24_leadingZeros_T_93[6] ? 6'h6 : _ans_24_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_185 = _ans_24_leadingZeros_T_93[5] ? 6'h5 : _ans_24_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_186 = _ans_24_leadingZeros_T_93[4] ? 6'h4 : _ans_24_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_187 = _ans_24_leadingZeros_T_93[3] ? 6'h3 : _ans_24_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_188 = _ans_24_leadingZeros_T_93[2] ? 6'h2 : _ans_24_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_leadingZeros_T_189 = _ans_24_leadingZeros_T_93[1] ? 6'h1 : _ans_24_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_24_leadingZeros = _ans_24_leadingZeros_T_93[0] ? 6'h0 : _ans_24_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_24_expRaw_T_1 = 6'h1f - ans_24_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_24_expRaw = ans_24_isZero ? 6'h0 : _ans_24_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_24_shiftAmt_T_2 = ans_24_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_24_shiftAmt = ans_24_expRaw > 6'h3 ? _ans_24_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_24_mantissaRaw_T = ans_24_absClipped >> ans_24_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_24_mantissaRaw = _ans_24_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_24_mantissa = ans_24_expRaw >= 6'h3 ? ans_24_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_24_expAdjusted = ans_24_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_24_exp_T_4 = ans_24_expAdjusted > 7'hf ? 4'hf : ans_24_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_24_exp = ans_24_isZero ? 4'h0 : _ans_24_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_24_fp8 = {ans_24_clippedX[31],ans_24_exp,ans_24_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_25 = {24'h0,linear_bias_25}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_25 = tempSum_25 + biasExtended_25; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_25_sign = sum32_25[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_25_absX_T = ~sum32_25; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_25_absX_T_2 = _ans_25_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_25_absX = ans_25_sign ? _ans_25_absX_T_2 : sum32_25; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_25_shiftedX_T_1 = _GEN_14432 - ans_25_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_25_shiftedX_T_3 = ans_25_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_25_shiftedX = ans_25_sign ? _ans_25_shiftedX_T_1 : _ans_25_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_25_scaledX_T_1 = ans_25_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_25_scaledX = _ans_25_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_25_clippedX_T_2 = ans_25_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_25_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_25_clippedX = ans_25_scaledX > 49'h1c0 ? 49'h1c0 : _ans_25_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_25_absClipped_T_1 = ~ans_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_25_absClipped_T_3 = _ans_25_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_25_absClipped = ans_25_clippedX[31] ? _ans_25_absClipped_T_3 : ans_25_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_25_isZero = ans_25_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_39989 = {{16'd0}, ans_25_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_4 = _GEN_39989 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_6 = {ans_25_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_8 = _ans_25_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_9 = _ans_25_leadingZeros_T_4 | _ans_25_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39990 = {{8'd0}, _ans_25_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_14 = _GEN_39990 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_16 = {_ans_25_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_18 = _ans_25_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_19 = _ans_25_leadingZeros_T_14 | _ans_25_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39991 = {{4'd0}, _ans_25_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_24 = _GEN_39991 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_26 = {_ans_25_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_28 = _ans_25_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_29 = _ans_25_leadingZeros_T_24 | _ans_25_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39992 = {{2'd0}, _ans_25_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_34 = _GEN_39992 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_36 = {_ans_25_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_38 = _ans_25_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_39 = _ans_25_leadingZeros_T_34 | _ans_25_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_39993 = {{1'd0}, _ans_25_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_44 = _GEN_39993 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_46 = {_ans_25_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_48 = _ans_25_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_25_leadingZeros_T_49 = _ans_25_leadingZeros_T_44 | _ans_25_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39994 = {{8'd0}, ans_25_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_55 = _GEN_39994 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_57 = {ans_25_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_59 = _ans_25_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_60 = _ans_25_leadingZeros_T_55 | _ans_25_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39995 = {{4'd0}, _ans_25_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_65 = _GEN_39995 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_67 = {_ans_25_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_69 = _ans_25_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_70 = _ans_25_leadingZeros_T_65 | _ans_25_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39996 = {{2'd0}, _ans_25_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_75 = _GEN_39996 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_77 = {_ans_25_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_79 = _ans_25_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_80 = _ans_25_leadingZeros_T_75 | _ans_25_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_39997 = {{1'd0}, _ans_25_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_85 = _GEN_39997 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_87 = {_ans_25_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_89 = _ans_25_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_25_leadingZeros_T_90 = _ans_25_leadingZeros_T_85 | _ans_25_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_25_leadingZeros_T_93 = {_ans_25_leadingZeros_T_49,_ans_25_leadingZeros_T_90,ans_25_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_25_leadingZeros_T_143 = _ans_25_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_144 = _ans_25_leadingZeros_T_93[46] ? 6'h2e : _ans_25_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_145 = _ans_25_leadingZeros_T_93[45] ? 6'h2d : _ans_25_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_146 = _ans_25_leadingZeros_T_93[44] ? 6'h2c : _ans_25_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_147 = _ans_25_leadingZeros_T_93[43] ? 6'h2b : _ans_25_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_148 = _ans_25_leadingZeros_T_93[42] ? 6'h2a : _ans_25_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_149 = _ans_25_leadingZeros_T_93[41] ? 6'h29 : _ans_25_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_150 = _ans_25_leadingZeros_T_93[40] ? 6'h28 : _ans_25_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_151 = _ans_25_leadingZeros_T_93[39] ? 6'h27 : _ans_25_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_152 = _ans_25_leadingZeros_T_93[38] ? 6'h26 : _ans_25_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_153 = _ans_25_leadingZeros_T_93[37] ? 6'h25 : _ans_25_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_154 = _ans_25_leadingZeros_T_93[36] ? 6'h24 : _ans_25_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_155 = _ans_25_leadingZeros_T_93[35] ? 6'h23 : _ans_25_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_156 = _ans_25_leadingZeros_T_93[34] ? 6'h22 : _ans_25_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_157 = _ans_25_leadingZeros_T_93[33] ? 6'h21 : _ans_25_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_158 = _ans_25_leadingZeros_T_93[32] ? 6'h20 : _ans_25_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_159 = _ans_25_leadingZeros_T_93[31] ? 6'h1f : _ans_25_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_160 = _ans_25_leadingZeros_T_93[30] ? 6'h1e : _ans_25_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_161 = _ans_25_leadingZeros_T_93[29] ? 6'h1d : _ans_25_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_162 = _ans_25_leadingZeros_T_93[28] ? 6'h1c : _ans_25_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_163 = _ans_25_leadingZeros_T_93[27] ? 6'h1b : _ans_25_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_164 = _ans_25_leadingZeros_T_93[26] ? 6'h1a : _ans_25_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_165 = _ans_25_leadingZeros_T_93[25] ? 6'h19 : _ans_25_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_166 = _ans_25_leadingZeros_T_93[24] ? 6'h18 : _ans_25_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_167 = _ans_25_leadingZeros_T_93[23] ? 6'h17 : _ans_25_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_168 = _ans_25_leadingZeros_T_93[22] ? 6'h16 : _ans_25_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_169 = _ans_25_leadingZeros_T_93[21] ? 6'h15 : _ans_25_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_170 = _ans_25_leadingZeros_T_93[20] ? 6'h14 : _ans_25_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_171 = _ans_25_leadingZeros_T_93[19] ? 6'h13 : _ans_25_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_172 = _ans_25_leadingZeros_T_93[18] ? 6'h12 : _ans_25_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_173 = _ans_25_leadingZeros_T_93[17] ? 6'h11 : _ans_25_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_174 = _ans_25_leadingZeros_T_93[16] ? 6'h10 : _ans_25_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_175 = _ans_25_leadingZeros_T_93[15] ? 6'hf : _ans_25_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_176 = _ans_25_leadingZeros_T_93[14] ? 6'he : _ans_25_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_177 = _ans_25_leadingZeros_T_93[13] ? 6'hd : _ans_25_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_178 = _ans_25_leadingZeros_T_93[12] ? 6'hc : _ans_25_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_179 = _ans_25_leadingZeros_T_93[11] ? 6'hb : _ans_25_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_180 = _ans_25_leadingZeros_T_93[10] ? 6'ha : _ans_25_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_181 = _ans_25_leadingZeros_T_93[9] ? 6'h9 : _ans_25_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_182 = _ans_25_leadingZeros_T_93[8] ? 6'h8 : _ans_25_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_183 = _ans_25_leadingZeros_T_93[7] ? 6'h7 : _ans_25_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_184 = _ans_25_leadingZeros_T_93[6] ? 6'h6 : _ans_25_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_185 = _ans_25_leadingZeros_T_93[5] ? 6'h5 : _ans_25_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_186 = _ans_25_leadingZeros_T_93[4] ? 6'h4 : _ans_25_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_187 = _ans_25_leadingZeros_T_93[3] ? 6'h3 : _ans_25_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_188 = _ans_25_leadingZeros_T_93[2] ? 6'h2 : _ans_25_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_leadingZeros_T_189 = _ans_25_leadingZeros_T_93[1] ? 6'h1 : _ans_25_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_25_leadingZeros = _ans_25_leadingZeros_T_93[0] ? 6'h0 : _ans_25_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_25_expRaw_T_1 = 6'h1f - ans_25_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_25_expRaw = ans_25_isZero ? 6'h0 : _ans_25_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_25_shiftAmt_T_2 = ans_25_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_25_shiftAmt = ans_25_expRaw > 6'h3 ? _ans_25_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_25_mantissaRaw_T = ans_25_absClipped >> ans_25_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_25_mantissaRaw = _ans_25_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_25_mantissa = ans_25_expRaw >= 6'h3 ? ans_25_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_25_expAdjusted = ans_25_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_25_exp_T_4 = ans_25_expAdjusted > 7'hf ? 4'hf : ans_25_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_25_exp = ans_25_isZero ? 4'h0 : _ans_25_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_25_fp8 = {ans_25_clippedX[31],ans_25_exp,ans_25_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_26 = {24'h0,linear_bias_26}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_26 = tempSum_26 + biasExtended_26; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_26_sign = sum32_26[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_26_absX_T = ~sum32_26; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_26_absX_T_2 = _ans_26_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_26_absX = ans_26_sign ? _ans_26_absX_T_2 : sum32_26; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_26_shiftedX_T_1 = _GEN_14432 - ans_26_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_26_shiftedX_T_3 = ans_26_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_26_shiftedX = ans_26_sign ? _ans_26_shiftedX_T_1 : _ans_26_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_26_scaledX_T_1 = ans_26_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_26_scaledX = _ans_26_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_26_clippedX_T_2 = ans_26_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_26_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_26_clippedX = ans_26_scaledX > 49'h1c0 ? 49'h1c0 : _ans_26_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_26_absClipped_T_1 = ~ans_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_26_absClipped_T_3 = _ans_26_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_26_absClipped = ans_26_clippedX[31] ? _ans_26_absClipped_T_3 : ans_26_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_26_isZero = ans_26_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40000 = {{16'd0}, ans_26_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_4 = _GEN_40000 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_6 = {ans_26_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_8 = _ans_26_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_9 = _ans_26_leadingZeros_T_4 | _ans_26_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40001 = {{8'd0}, _ans_26_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_14 = _GEN_40001 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_16 = {_ans_26_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_18 = _ans_26_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_19 = _ans_26_leadingZeros_T_14 | _ans_26_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40002 = {{4'd0}, _ans_26_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_24 = _GEN_40002 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_26 = {_ans_26_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_28 = _ans_26_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_29 = _ans_26_leadingZeros_T_24 | _ans_26_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40003 = {{2'd0}, _ans_26_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_34 = _GEN_40003 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_36 = {_ans_26_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_38 = _ans_26_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_39 = _ans_26_leadingZeros_T_34 | _ans_26_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40004 = {{1'd0}, _ans_26_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_44 = _GEN_40004 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_46 = {_ans_26_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_48 = _ans_26_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_26_leadingZeros_T_49 = _ans_26_leadingZeros_T_44 | _ans_26_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40005 = {{8'd0}, ans_26_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_55 = _GEN_40005 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_57 = {ans_26_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_59 = _ans_26_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_60 = _ans_26_leadingZeros_T_55 | _ans_26_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40006 = {{4'd0}, _ans_26_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_65 = _GEN_40006 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_67 = {_ans_26_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_69 = _ans_26_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_70 = _ans_26_leadingZeros_T_65 | _ans_26_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40007 = {{2'd0}, _ans_26_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_75 = _GEN_40007 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_77 = {_ans_26_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_79 = _ans_26_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_80 = _ans_26_leadingZeros_T_75 | _ans_26_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40008 = {{1'd0}, _ans_26_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_85 = _GEN_40008 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_87 = {_ans_26_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_89 = _ans_26_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_26_leadingZeros_T_90 = _ans_26_leadingZeros_T_85 | _ans_26_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_26_leadingZeros_T_93 = {_ans_26_leadingZeros_T_49,_ans_26_leadingZeros_T_90,ans_26_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_26_leadingZeros_T_143 = _ans_26_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_144 = _ans_26_leadingZeros_T_93[46] ? 6'h2e : _ans_26_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_145 = _ans_26_leadingZeros_T_93[45] ? 6'h2d : _ans_26_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_146 = _ans_26_leadingZeros_T_93[44] ? 6'h2c : _ans_26_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_147 = _ans_26_leadingZeros_T_93[43] ? 6'h2b : _ans_26_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_148 = _ans_26_leadingZeros_T_93[42] ? 6'h2a : _ans_26_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_149 = _ans_26_leadingZeros_T_93[41] ? 6'h29 : _ans_26_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_150 = _ans_26_leadingZeros_T_93[40] ? 6'h28 : _ans_26_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_151 = _ans_26_leadingZeros_T_93[39] ? 6'h27 : _ans_26_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_152 = _ans_26_leadingZeros_T_93[38] ? 6'h26 : _ans_26_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_153 = _ans_26_leadingZeros_T_93[37] ? 6'h25 : _ans_26_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_154 = _ans_26_leadingZeros_T_93[36] ? 6'h24 : _ans_26_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_155 = _ans_26_leadingZeros_T_93[35] ? 6'h23 : _ans_26_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_156 = _ans_26_leadingZeros_T_93[34] ? 6'h22 : _ans_26_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_157 = _ans_26_leadingZeros_T_93[33] ? 6'h21 : _ans_26_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_158 = _ans_26_leadingZeros_T_93[32] ? 6'h20 : _ans_26_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_159 = _ans_26_leadingZeros_T_93[31] ? 6'h1f : _ans_26_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_160 = _ans_26_leadingZeros_T_93[30] ? 6'h1e : _ans_26_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_161 = _ans_26_leadingZeros_T_93[29] ? 6'h1d : _ans_26_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_162 = _ans_26_leadingZeros_T_93[28] ? 6'h1c : _ans_26_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_163 = _ans_26_leadingZeros_T_93[27] ? 6'h1b : _ans_26_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_164 = _ans_26_leadingZeros_T_93[26] ? 6'h1a : _ans_26_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_165 = _ans_26_leadingZeros_T_93[25] ? 6'h19 : _ans_26_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_166 = _ans_26_leadingZeros_T_93[24] ? 6'h18 : _ans_26_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_167 = _ans_26_leadingZeros_T_93[23] ? 6'h17 : _ans_26_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_168 = _ans_26_leadingZeros_T_93[22] ? 6'h16 : _ans_26_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_169 = _ans_26_leadingZeros_T_93[21] ? 6'h15 : _ans_26_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_170 = _ans_26_leadingZeros_T_93[20] ? 6'h14 : _ans_26_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_171 = _ans_26_leadingZeros_T_93[19] ? 6'h13 : _ans_26_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_172 = _ans_26_leadingZeros_T_93[18] ? 6'h12 : _ans_26_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_173 = _ans_26_leadingZeros_T_93[17] ? 6'h11 : _ans_26_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_174 = _ans_26_leadingZeros_T_93[16] ? 6'h10 : _ans_26_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_175 = _ans_26_leadingZeros_T_93[15] ? 6'hf : _ans_26_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_176 = _ans_26_leadingZeros_T_93[14] ? 6'he : _ans_26_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_177 = _ans_26_leadingZeros_T_93[13] ? 6'hd : _ans_26_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_178 = _ans_26_leadingZeros_T_93[12] ? 6'hc : _ans_26_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_179 = _ans_26_leadingZeros_T_93[11] ? 6'hb : _ans_26_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_180 = _ans_26_leadingZeros_T_93[10] ? 6'ha : _ans_26_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_181 = _ans_26_leadingZeros_T_93[9] ? 6'h9 : _ans_26_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_182 = _ans_26_leadingZeros_T_93[8] ? 6'h8 : _ans_26_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_183 = _ans_26_leadingZeros_T_93[7] ? 6'h7 : _ans_26_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_184 = _ans_26_leadingZeros_T_93[6] ? 6'h6 : _ans_26_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_185 = _ans_26_leadingZeros_T_93[5] ? 6'h5 : _ans_26_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_186 = _ans_26_leadingZeros_T_93[4] ? 6'h4 : _ans_26_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_187 = _ans_26_leadingZeros_T_93[3] ? 6'h3 : _ans_26_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_188 = _ans_26_leadingZeros_T_93[2] ? 6'h2 : _ans_26_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_leadingZeros_T_189 = _ans_26_leadingZeros_T_93[1] ? 6'h1 : _ans_26_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_26_leadingZeros = _ans_26_leadingZeros_T_93[0] ? 6'h0 : _ans_26_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_26_expRaw_T_1 = 6'h1f - ans_26_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_26_expRaw = ans_26_isZero ? 6'h0 : _ans_26_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_26_shiftAmt_T_2 = ans_26_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_26_shiftAmt = ans_26_expRaw > 6'h3 ? _ans_26_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_26_mantissaRaw_T = ans_26_absClipped >> ans_26_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_26_mantissaRaw = _ans_26_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_26_mantissa = ans_26_expRaw >= 6'h3 ? ans_26_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_26_expAdjusted = ans_26_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_26_exp_T_4 = ans_26_expAdjusted > 7'hf ? 4'hf : ans_26_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_26_exp = ans_26_isZero ? 4'h0 : _ans_26_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_26_fp8 = {ans_26_clippedX[31],ans_26_exp,ans_26_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_27 = {24'h0,linear_bias_27}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_27 = tempSum_27 + biasExtended_27; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_27_sign = sum32_27[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_27_absX_T = ~sum32_27; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_27_absX_T_2 = _ans_27_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_27_absX = ans_27_sign ? _ans_27_absX_T_2 : sum32_27; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_27_shiftedX_T_1 = _GEN_14432 - ans_27_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_27_shiftedX_T_3 = ans_27_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_27_shiftedX = ans_27_sign ? _ans_27_shiftedX_T_1 : _ans_27_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_27_scaledX_T_1 = ans_27_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_27_scaledX = _ans_27_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_27_clippedX_T_2 = ans_27_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_27_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_27_clippedX = ans_27_scaledX > 49'h1c0 ? 49'h1c0 : _ans_27_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_27_absClipped_T_1 = ~ans_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_27_absClipped_T_3 = _ans_27_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_27_absClipped = ans_27_clippedX[31] ? _ans_27_absClipped_T_3 : ans_27_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_27_isZero = ans_27_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40011 = {{16'd0}, ans_27_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_4 = _GEN_40011 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_6 = {ans_27_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_8 = _ans_27_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_9 = _ans_27_leadingZeros_T_4 | _ans_27_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40012 = {{8'd0}, _ans_27_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_14 = _GEN_40012 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_16 = {_ans_27_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_18 = _ans_27_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_19 = _ans_27_leadingZeros_T_14 | _ans_27_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40013 = {{4'd0}, _ans_27_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_24 = _GEN_40013 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_26 = {_ans_27_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_28 = _ans_27_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_29 = _ans_27_leadingZeros_T_24 | _ans_27_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40014 = {{2'd0}, _ans_27_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_34 = _GEN_40014 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_36 = {_ans_27_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_38 = _ans_27_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_39 = _ans_27_leadingZeros_T_34 | _ans_27_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40015 = {{1'd0}, _ans_27_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_44 = _GEN_40015 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_46 = {_ans_27_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_48 = _ans_27_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_27_leadingZeros_T_49 = _ans_27_leadingZeros_T_44 | _ans_27_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40016 = {{8'd0}, ans_27_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_55 = _GEN_40016 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_57 = {ans_27_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_59 = _ans_27_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_60 = _ans_27_leadingZeros_T_55 | _ans_27_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40017 = {{4'd0}, _ans_27_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_65 = _GEN_40017 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_67 = {_ans_27_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_69 = _ans_27_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_70 = _ans_27_leadingZeros_T_65 | _ans_27_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40018 = {{2'd0}, _ans_27_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_75 = _GEN_40018 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_77 = {_ans_27_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_79 = _ans_27_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_80 = _ans_27_leadingZeros_T_75 | _ans_27_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40019 = {{1'd0}, _ans_27_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_85 = _GEN_40019 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_87 = {_ans_27_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_89 = _ans_27_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_27_leadingZeros_T_90 = _ans_27_leadingZeros_T_85 | _ans_27_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_27_leadingZeros_T_93 = {_ans_27_leadingZeros_T_49,_ans_27_leadingZeros_T_90,ans_27_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_27_leadingZeros_T_143 = _ans_27_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_144 = _ans_27_leadingZeros_T_93[46] ? 6'h2e : _ans_27_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_145 = _ans_27_leadingZeros_T_93[45] ? 6'h2d : _ans_27_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_146 = _ans_27_leadingZeros_T_93[44] ? 6'h2c : _ans_27_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_147 = _ans_27_leadingZeros_T_93[43] ? 6'h2b : _ans_27_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_148 = _ans_27_leadingZeros_T_93[42] ? 6'h2a : _ans_27_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_149 = _ans_27_leadingZeros_T_93[41] ? 6'h29 : _ans_27_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_150 = _ans_27_leadingZeros_T_93[40] ? 6'h28 : _ans_27_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_151 = _ans_27_leadingZeros_T_93[39] ? 6'h27 : _ans_27_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_152 = _ans_27_leadingZeros_T_93[38] ? 6'h26 : _ans_27_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_153 = _ans_27_leadingZeros_T_93[37] ? 6'h25 : _ans_27_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_154 = _ans_27_leadingZeros_T_93[36] ? 6'h24 : _ans_27_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_155 = _ans_27_leadingZeros_T_93[35] ? 6'h23 : _ans_27_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_156 = _ans_27_leadingZeros_T_93[34] ? 6'h22 : _ans_27_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_157 = _ans_27_leadingZeros_T_93[33] ? 6'h21 : _ans_27_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_158 = _ans_27_leadingZeros_T_93[32] ? 6'h20 : _ans_27_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_159 = _ans_27_leadingZeros_T_93[31] ? 6'h1f : _ans_27_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_160 = _ans_27_leadingZeros_T_93[30] ? 6'h1e : _ans_27_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_161 = _ans_27_leadingZeros_T_93[29] ? 6'h1d : _ans_27_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_162 = _ans_27_leadingZeros_T_93[28] ? 6'h1c : _ans_27_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_163 = _ans_27_leadingZeros_T_93[27] ? 6'h1b : _ans_27_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_164 = _ans_27_leadingZeros_T_93[26] ? 6'h1a : _ans_27_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_165 = _ans_27_leadingZeros_T_93[25] ? 6'h19 : _ans_27_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_166 = _ans_27_leadingZeros_T_93[24] ? 6'h18 : _ans_27_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_167 = _ans_27_leadingZeros_T_93[23] ? 6'h17 : _ans_27_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_168 = _ans_27_leadingZeros_T_93[22] ? 6'h16 : _ans_27_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_169 = _ans_27_leadingZeros_T_93[21] ? 6'h15 : _ans_27_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_170 = _ans_27_leadingZeros_T_93[20] ? 6'h14 : _ans_27_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_171 = _ans_27_leadingZeros_T_93[19] ? 6'h13 : _ans_27_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_172 = _ans_27_leadingZeros_T_93[18] ? 6'h12 : _ans_27_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_173 = _ans_27_leadingZeros_T_93[17] ? 6'h11 : _ans_27_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_174 = _ans_27_leadingZeros_T_93[16] ? 6'h10 : _ans_27_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_175 = _ans_27_leadingZeros_T_93[15] ? 6'hf : _ans_27_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_176 = _ans_27_leadingZeros_T_93[14] ? 6'he : _ans_27_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_177 = _ans_27_leadingZeros_T_93[13] ? 6'hd : _ans_27_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_178 = _ans_27_leadingZeros_T_93[12] ? 6'hc : _ans_27_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_179 = _ans_27_leadingZeros_T_93[11] ? 6'hb : _ans_27_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_180 = _ans_27_leadingZeros_T_93[10] ? 6'ha : _ans_27_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_181 = _ans_27_leadingZeros_T_93[9] ? 6'h9 : _ans_27_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_182 = _ans_27_leadingZeros_T_93[8] ? 6'h8 : _ans_27_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_183 = _ans_27_leadingZeros_T_93[7] ? 6'h7 : _ans_27_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_184 = _ans_27_leadingZeros_T_93[6] ? 6'h6 : _ans_27_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_185 = _ans_27_leadingZeros_T_93[5] ? 6'h5 : _ans_27_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_186 = _ans_27_leadingZeros_T_93[4] ? 6'h4 : _ans_27_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_187 = _ans_27_leadingZeros_T_93[3] ? 6'h3 : _ans_27_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_188 = _ans_27_leadingZeros_T_93[2] ? 6'h2 : _ans_27_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_leadingZeros_T_189 = _ans_27_leadingZeros_T_93[1] ? 6'h1 : _ans_27_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_27_leadingZeros = _ans_27_leadingZeros_T_93[0] ? 6'h0 : _ans_27_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_27_expRaw_T_1 = 6'h1f - ans_27_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_27_expRaw = ans_27_isZero ? 6'h0 : _ans_27_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_27_shiftAmt_T_2 = ans_27_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_27_shiftAmt = ans_27_expRaw > 6'h3 ? _ans_27_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_27_mantissaRaw_T = ans_27_absClipped >> ans_27_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_27_mantissaRaw = _ans_27_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_27_mantissa = ans_27_expRaw >= 6'h3 ? ans_27_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_27_expAdjusted = ans_27_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_27_exp_T_4 = ans_27_expAdjusted > 7'hf ? 4'hf : ans_27_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_27_exp = ans_27_isZero ? 4'h0 : _ans_27_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_27_fp8 = {ans_27_clippedX[31],ans_27_exp,ans_27_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_28 = {24'h0,linear_bias_28}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_28 = tempSum_28 + biasExtended_28; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_28_sign = sum32_28[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_28_absX_T = ~sum32_28; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_28_absX_T_2 = _ans_28_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_28_absX = ans_28_sign ? _ans_28_absX_T_2 : sum32_28; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_28_shiftedX_T_1 = _GEN_14432 - ans_28_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_28_shiftedX_T_3 = ans_28_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_28_shiftedX = ans_28_sign ? _ans_28_shiftedX_T_1 : _ans_28_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_28_scaledX_T_1 = ans_28_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_28_scaledX = _ans_28_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_28_clippedX_T_2 = ans_28_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_28_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_28_clippedX = ans_28_scaledX > 49'h1c0 ? 49'h1c0 : _ans_28_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_28_absClipped_T_1 = ~ans_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_28_absClipped_T_3 = _ans_28_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_28_absClipped = ans_28_clippedX[31] ? _ans_28_absClipped_T_3 : ans_28_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_28_isZero = ans_28_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40022 = {{16'd0}, ans_28_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_4 = _GEN_40022 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_6 = {ans_28_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_8 = _ans_28_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_9 = _ans_28_leadingZeros_T_4 | _ans_28_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40023 = {{8'd0}, _ans_28_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_14 = _GEN_40023 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_16 = {_ans_28_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_18 = _ans_28_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_19 = _ans_28_leadingZeros_T_14 | _ans_28_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40024 = {{4'd0}, _ans_28_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_24 = _GEN_40024 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_26 = {_ans_28_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_28 = _ans_28_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_29 = _ans_28_leadingZeros_T_24 | _ans_28_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40025 = {{2'd0}, _ans_28_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_34 = _GEN_40025 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_36 = {_ans_28_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_38 = _ans_28_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_39 = _ans_28_leadingZeros_T_34 | _ans_28_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40026 = {{1'd0}, _ans_28_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_44 = _GEN_40026 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_46 = {_ans_28_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_48 = _ans_28_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_28_leadingZeros_T_49 = _ans_28_leadingZeros_T_44 | _ans_28_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40027 = {{8'd0}, ans_28_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_55 = _GEN_40027 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_57 = {ans_28_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_59 = _ans_28_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_60 = _ans_28_leadingZeros_T_55 | _ans_28_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40028 = {{4'd0}, _ans_28_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_65 = _GEN_40028 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_67 = {_ans_28_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_69 = _ans_28_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_70 = _ans_28_leadingZeros_T_65 | _ans_28_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40029 = {{2'd0}, _ans_28_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_75 = _GEN_40029 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_77 = {_ans_28_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_79 = _ans_28_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_80 = _ans_28_leadingZeros_T_75 | _ans_28_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40030 = {{1'd0}, _ans_28_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_85 = _GEN_40030 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_87 = {_ans_28_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_89 = _ans_28_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_28_leadingZeros_T_90 = _ans_28_leadingZeros_T_85 | _ans_28_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_28_leadingZeros_T_93 = {_ans_28_leadingZeros_T_49,_ans_28_leadingZeros_T_90,ans_28_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_28_leadingZeros_T_143 = _ans_28_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_144 = _ans_28_leadingZeros_T_93[46] ? 6'h2e : _ans_28_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_145 = _ans_28_leadingZeros_T_93[45] ? 6'h2d : _ans_28_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_146 = _ans_28_leadingZeros_T_93[44] ? 6'h2c : _ans_28_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_147 = _ans_28_leadingZeros_T_93[43] ? 6'h2b : _ans_28_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_148 = _ans_28_leadingZeros_T_93[42] ? 6'h2a : _ans_28_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_149 = _ans_28_leadingZeros_T_93[41] ? 6'h29 : _ans_28_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_150 = _ans_28_leadingZeros_T_93[40] ? 6'h28 : _ans_28_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_151 = _ans_28_leadingZeros_T_93[39] ? 6'h27 : _ans_28_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_152 = _ans_28_leadingZeros_T_93[38] ? 6'h26 : _ans_28_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_153 = _ans_28_leadingZeros_T_93[37] ? 6'h25 : _ans_28_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_154 = _ans_28_leadingZeros_T_93[36] ? 6'h24 : _ans_28_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_155 = _ans_28_leadingZeros_T_93[35] ? 6'h23 : _ans_28_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_156 = _ans_28_leadingZeros_T_93[34] ? 6'h22 : _ans_28_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_157 = _ans_28_leadingZeros_T_93[33] ? 6'h21 : _ans_28_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_158 = _ans_28_leadingZeros_T_93[32] ? 6'h20 : _ans_28_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_159 = _ans_28_leadingZeros_T_93[31] ? 6'h1f : _ans_28_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_160 = _ans_28_leadingZeros_T_93[30] ? 6'h1e : _ans_28_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_161 = _ans_28_leadingZeros_T_93[29] ? 6'h1d : _ans_28_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_162 = _ans_28_leadingZeros_T_93[28] ? 6'h1c : _ans_28_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_163 = _ans_28_leadingZeros_T_93[27] ? 6'h1b : _ans_28_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_164 = _ans_28_leadingZeros_T_93[26] ? 6'h1a : _ans_28_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_165 = _ans_28_leadingZeros_T_93[25] ? 6'h19 : _ans_28_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_166 = _ans_28_leadingZeros_T_93[24] ? 6'h18 : _ans_28_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_167 = _ans_28_leadingZeros_T_93[23] ? 6'h17 : _ans_28_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_168 = _ans_28_leadingZeros_T_93[22] ? 6'h16 : _ans_28_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_169 = _ans_28_leadingZeros_T_93[21] ? 6'h15 : _ans_28_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_170 = _ans_28_leadingZeros_T_93[20] ? 6'h14 : _ans_28_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_171 = _ans_28_leadingZeros_T_93[19] ? 6'h13 : _ans_28_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_172 = _ans_28_leadingZeros_T_93[18] ? 6'h12 : _ans_28_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_173 = _ans_28_leadingZeros_T_93[17] ? 6'h11 : _ans_28_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_174 = _ans_28_leadingZeros_T_93[16] ? 6'h10 : _ans_28_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_175 = _ans_28_leadingZeros_T_93[15] ? 6'hf : _ans_28_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_176 = _ans_28_leadingZeros_T_93[14] ? 6'he : _ans_28_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_177 = _ans_28_leadingZeros_T_93[13] ? 6'hd : _ans_28_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_178 = _ans_28_leadingZeros_T_93[12] ? 6'hc : _ans_28_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_179 = _ans_28_leadingZeros_T_93[11] ? 6'hb : _ans_28_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_180 = _ans_28_leadingZeros_T_93[10] ? 6'ha : _ans_28_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_181 = _ans_28_leadingZeros_T_93[9] ? 6'h9 : _ans_28_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_182 = _ans_28_leadingZeros_T_93[8] ? 6'h8 : _ans_28_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_183 = _ans_28_leadingZeros_T_93[7] ? 6'h7 : _ans_28_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_184 = _ans_28_leadingZeros_T_93[6] ? 6'h6 : _ans_28_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_185 = _ans_28_leadingZeros_T_93[5] ? 6'h5 : _ans_28_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_186 = _ans_28_leadingZeros_T_93[4] ? 6'h4 : _ans_28_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_187 = _ans_28_leadingZeros_T_93[3] ? 6'h3 : _ans_28_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_188 = _ans_28_leadingZeros_T_93[2] ? 6'h2 : _ans_28_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_leadingZeros_T_189 = _ans_28_leadingZeros_T_93[1] ? 6'h1 : _ans_28_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_28_leadingZeros = _ans_28_leadingZeros_T_93[0] ? 6'h0 : _ans_28_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_28_expRaw_T_1 = 6'h1f - ans_28_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_28_expRaw = ans_28_isZero ? 6'h0 : _ans_28_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_28_shiftAmt_T_2 = ans_28_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_28_shiftAmt = ans_28_expRaw > 6'h3 ? _ans_28_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_28_mantissaRaw_T = ans_28_absClipped >> ans_28_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_28_mantissaRaw = _ans_28_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_28_mantissa = ans_28_expRaw >= 6'h3 ? ans_28_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_28_expAdjusted = ans_28_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_28_exp_T_4 = ans_28_expAdjusted > 7'hf ? 4'hf : ans_28_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_28_exp = ans_28_isZero ? 4'h0 : _ans_28_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_28_fp8 = {ans_28_clippedX[31],ans_28_exp,ans_28_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_29 = {24'h0,linear_bias_29}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_29 = tempSum_29 + biasExtended_29; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_29_sign = sum32_29[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_29_absX_T = ~sum32_29; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_29_absX_T_2 = _ans_29_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_29_absX = ans_29_sign ? _ans_29_absX_T_2 : sum32_29; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_29_shiftedX_T_1 = _GEN_14432 - ans_29_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_29_shiftedX_T_3 = ans_29_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_29_shiftedX = ans_29_sign ? _ans_29_shiftedX_T_1 : _ans_29_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_29_scaledX_T_1 = ans_29_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_29_scaledX = _ans_29_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_29_clippedX_T_2 = ans_29_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_29_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_29_clippedX = ans_29_scaledX > 49'h1c0 ? 49'h1c0 : _ans_29_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_29_absClipped_T_1 = ~ans_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_29_absClipped_T_3 = _ans_29_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_29_absClipped = ans_29_clippedX[31] ? _ans_29_absClipped_T_3 : ans_29_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_29_isZero = ans_29_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40033 = {{16'd0}, ans_29_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_4 = _GEN_40033 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_6 = {ans_29_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_8 = _ans_29_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_9 = _ans_29_leadingZeros_T_4 | _ans_29_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40034 = {{8'd0}, _ans_29_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_14 = _GEN_40034 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_16 = {_ans_29_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_18 = _ans_29_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_19 = _ans_29_leadingZeros_T_14 | _ans_29_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40035 = {{4'd0}, _ans_29_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_24 = _GEN_40035 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_26 = {_ans_29_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_28 = _ans_29_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_29 = _ans_29_leadingZeros_T_24 | _ans_29_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40036 = {{2'd0}, _ans_29_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_34 = _GEN_40036 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_36 = {_ans_29_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_38 = _ans_29_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_39 = _ans_29_leadingZeros_T_34 | _ans_29_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40037 = {{1'd0}, _ans_29_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_44 = _GEN_40037 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_46 = {_ans_29_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_48 = _ans_29_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_29_leadingZeros_T_49 = _ans_29_leadingZeros_T_44 | _ans_29_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40038 = {{8'd0}, ans_29_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_55 = _GEN_40038 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_57 = {ans_29_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_59 = _ans_29_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_60 = _ans_29_leadingZeros_T_55 | _ans_29_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40039 = {{4'd0}, _ans_29_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_65 = _GEN_40039 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_67 = {_ans_29_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_69 = _ans_29_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_70 = _ans_29_leadingZeros_T_65 | _ans_29_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40040 = {{2'd0}, _ans_29_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_75 = _GEN_40040 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_77 = {_ans_29_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_79 = _ans_29_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_80 = _ans_29_leadingZeros_T_75 | _ans_29_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40041 = {{1'd0}, _ans_29_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_85 = _GEN_40041 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_87 = {_ans_29_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_89 = _ans_29_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_29_leadingZeros_T_90 = _ans_29_leadingZeros_T_85 | _ans_29_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_29_leadingZeros_T_93 = {_ans_29_leadingZeros_T_49,_ans_29_leadingZeros_T_90,ans_29_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_29_leadingZeros_T_143 = _ans_29_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_144 = _ans_29_leadingZeros_T_93[46] ? 6'h2e : _ans_29_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_145 = _ans_29_leadingZeros_T_93[45] ? 6'h2d : _ans_29_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_146 = _ans_29_leadingZeros_T_93[44] ? 6'h2c : _ans_29_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_147 = _ans_29_leadingZeros_T_93[43] ? 6'h2b : _ans_29_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_148 = _ans_29_leadingZeros_T_93[42] ? 6'h2a : _ans_29_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_149 = _ans_29_leadingZeros_T_93[41] ? 6'h29 : _ans_29_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_150 = _ans_29_leadingZeros_T_93[40] ? 6'h28 : _ans_29_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_151 = _ans_29_leadingZeros_T_93[39] ? 6'h27 : _ans_29_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_152 = _ans_29_leadingZeros_T_93[38] ? 6'h26 : _ans_29_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_153 = _ans_29_leadingZeros_T_93[37] ? 6'h25 : _ans_29_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_154 = _ans_29_leadingZeros_T_93[36] ? 6'h24 : _ans_29_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_155 = _ans_29_leadingZeros_T_93[35] ? 6'h23 : _ans_29_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_156 = _ans_29_leadingZeros_T_93[34] ? 6'h22 : _ans_29_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_157 = _ans_29_leadingZeros_T_93[33] ? 6'h21 : _ans_29_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_158 = _ans_29_leadingZeros_T_93[32] ? 6'h20 : _ans_29_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_159 = _ans_29_leadingZeros_T_93[31] ? 6'h1f : _ans_29_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_160 = _ans_29_leadingZeros_T_93[30] ? 6'h1e : _ans_29_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_161 = _ans_29_leadingZeros_T_93[29] ? 6'h1d : _ans_29_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_162 = _ans_29_leadingZeros_T_93[28] ? 6'h1c : _ans_29_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_163 = _ans_29_leadingZeros_T_93[27] ? 6'h1b : _ans_29_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_164 = _ans_29_leadingZeros_T_93[26] ? 6'h1a : _ans_29_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_165 = _ans_29_leadingZeros_T_93[25] ? 6'h19 : _ans_29_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_166 = _ans_29_leadingZeros_T_93[24] ? 6'h18 : _ans_29_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_167 = _ans_29_leadingZeros_T_93[23] ? 6'h17 : _ans_29_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_168 = _ans_29_leadingZeros_T_93[22] ? 6'h16 : _ans_29_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_169 = _ans_29_leadingZeros_T_93[21] ? 6'h15 : _ans_29_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_170 = _ans_29_leadingZeros_T_93[20] ? 6'h14 : _ans_29_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_171 = _ans_29_leadingZeros_T_93[19] ? 6'h13 : _ans_29_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_172 = _ans_29_leadingZeros_T_93[18] ? 6'h12 : _ans_29_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_173 = _ans_29_leadingZeros_T_93[17] ? 6'h11 : _ans_29_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_174 = _ans_29_leadingZeros_T_93[16] ? 6'h10 : _ans_29_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_175 = _ans_29_leadingZeros_T_93[15] ? 6'hf : _ans_29_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_176 = _ans_29_leadingZeros_T_93[14] ? 6'he : _ans_29_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_177 = _ans_29_leadingZeros_T_93[13] ? 6'hd : _ans_29_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_178 = _ans_29_leadingZeros_T_93[12] ? 6'hc : _ans_29_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_179 = _ans_29_leadingZeros_T_93[11] ? 6'hb : _ans_29_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_180 = _ans_29_leadingZeros_T_93[10] ? 6'ha : _ans_29_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_181 = _ans_29_leadingZeros_T_93[9] ? 6'h9 : _ans_29_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_182 = _ans_29_leadingZeros_T_93[8] ? 6'h8 : _ans_29_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_183 = _ans_29_leadingZeros_T_93[7] ? 6'h7 : _ans_29_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_184 = _ans_29_leadingZeros_T_93[6] ? 6'h6 : _ans_29_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_185 = _ans_29_leadingZeros_T_93[5] ? 6'h5 : _ans_29_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_186 = _ans_29_leadingZeros_T_93[4] ? 6'h4 : _ans_29_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_187 = _ans_29_leadingZeros_T_93[3] ? 6'h3 : _ans_29_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_188 = _ans_29_leadingZeros_T_93[2] ? 6'h2 : _ans_29_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_leadingZeros_T_189 = _ans_29_leadingZeros_T_93[1] ? 6'h1 : _ans_29_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_29_leadingZeros = _ans_29_leadingZeros_T_93[0] ? 6'h0 : _ans_29_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_29_expRaw_T_1 = 6'h1f - ans_29_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_29_expRaw = ans_29_isZero ? 6'h0 : _ans_29_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_29_shiftAmt_T_2 = ans_29_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_29_shiftAmt = ans_29_expRaw > 6'h3 ? _ans_29_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_29_mantissaRaw_T = ans_29_absClipped >> ans_29_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_29_mantissaRaw = _ans_29_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_29_mantissa = ans_29_expRaw >= 6'h3 ? ans_29_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_29_expAdjusted = ans_29_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_29_exp_T_4 = ans_29_expAdjusted > 7'hf ? 4'hf : ans_29_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_29_exp = ans_29_isZero ? 4'h0 : _ans_29_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_29_fp8 = {ans_29_clippedX[31],ans_29_exp,ans_29_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_30 = {24'h0,linear_bias_30}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_30 = tempSum_30 + biasExtended_30; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_30_sign = sum32_30[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_30_absX_T = ~sum32_30; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_30_absX_T_2 = _ans_30_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_30_absX = ans_30_sign ? _ans_30_absX_T_2 : sum32_30; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_30_shiftedX_T_1 = _GEN_14432 - ans_30_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_30_shiftedX_T_3 = ans_30_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_30_shiftedX = ans_30_sign ? _ans_30_shiftedX_T_1 : _ans_30_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_30_scaledX_T_1 = ans_30_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_30_scaledX = _ans_30_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_30_clippedX_T_2 = ans_30_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_30_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_30_clippedX = ans_30_scaledX > 49'h1c0 ? 49'h1c0 : _ans_30_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_30_absClipped_T_1 = ~ans_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_30_absClipped_T_3 = _ans_30_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_30_absClipped = ans_30_clippedX[31] ? _ans_30_absClipped_T_3 : ans_30_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_30_isZero = ans_30_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40044 = {{16'd0}, ans_30_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_4 = _GEN_40044 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_6 = {ans_30_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_8 = _ans_30_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_9 = _ans_30_leadingZeros_T_4 | _ans_30_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40045 = {{8'd0}, _ans_30_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_14 = _GEN_40045 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_16 = {_ans_30_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_18 = _ans_30_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_19 = _ans_30_leadingZeros_T_14 | _ans_30_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40046 = {{4'd0}, _ans_30_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_24 = _GEN_40046 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_26 = {_ans_30_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_28 = _ans_30_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_29 = _ans_30_leadingZeros_T_24 | _ans_30_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40047 = {{2'd0}, _ans_30_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_34 = _GEN_40047 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_36 = {_ans_30_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_38 = _ans_30_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_39 = _ans_30_leadingZeros_T_34 | _ans_30_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40048 = {{1'd0}, _ans_30_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_44 = _GEN_40048 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_46 = {_ans_30_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_48 = _ans_30_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_30_leadingZeros_T_49 = _ans_30_leadingZeros_T_44 | _ans_30_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40049 = {{8'd0}, ans_30_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_55 = _GEN_40049 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_57 = {ans_30_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_59 = _ans_30_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_60 = _ans_30_leadingZeros_T_55 | _ans_30_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40050 = {{4'd0}, _ans_30_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_65 = _GEN_40050 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_67 = {_ans_30_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_69 = _ans_30_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_70 = _ans_30_leadingZeros_T_65 | _ans_30_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40051 = {{2'd0}, _ans_30_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_75 = _GEN_40051 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_77 = {_ans_30_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_79 = _ans_30_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_80 = _ans_30_leadingZeros_T_75 | _ans_30_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40052 = {{1'd0}, _ans_30_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_85 = _GEN_40052 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_87 = {_ans_30_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_89 = _ans_30_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_30_leadingZeros_T_90 = _ans_30_leadingZeros_T_85 | _ans_30_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_30_leadingZeros_T_93 = {_ans_30_leadingZeros_T_49,_ans_30_leadingZeros_T_90,ans_30_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_30_leadingZeros_T_143 = _ans_30_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_144 = _ans_30_leadingZeros_T_93[46] ? 6'h2e : _ans_30_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_145 = _ans_30_leadingZeros_T_93[45] ? 6'h2d : _ans_30_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_146 = _ans_30_leadingZeros_T_93[44] ? 6'h2c : _ans_30_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_147 = _ans_30_leadingZeros_T_93[43] ? 6'h2b : _ans_30_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_148 = _ans_30_leadingZeros_T_93[42] ? 6'h2a : _ans_30_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_149 = _ans_30_leadingZeros_T_93[41] ? 6'h29 : _ans_30_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_150 = _ans_30_leadingZeros_T_93[40] ? 6'h28 : _ans_30_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_151 = _ans_30_leadingZeros_T_93[39] ? 6'h27 : _ans_30_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_152 = _ans_30_leadingZeros_T_93[38] ? 6'h26 : _ans_30_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_153 = _ans_30_leadingZeros_T_93[37] ? 6'h25 : _ans_30_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_154 = _ans_30_leadingZeros_T_93[36] ? 6'h24 : _ans_30_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_155 = _ans_30_leadingZeros_T_93[35] ? 6'h23 : _ans_30_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_156 = _ans_30_leadingZeros_T_93[34] ? 6'h22 : _ans_30_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_157 = _ans_30_leadingZeros_T_93[33] ? 6'h21 : _ans_30_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_158 = _ans_30_leadingZeros_T_93[32] ? 6'h20 : _ans_30_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_159 = _ans_30_leadingZeros_T_93[31] ? 6'h1f : _ans_30_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_160 = _ans_30_leadingZeros_T_93[30] ? 6'h1e : _ans_30_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_161 = _ans_30_leadingZeros_T_93[29] ? 6'h1d : _ans_30_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_162 = _ans_30_leadingZeros_T_93[28] ? 6'h1c : _ans_30_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_163 = _ans_30_leadingZeros_T_93[27] ? 6'h1b : _ans_30_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_164 = _ans_30_leadingZeros_T_93[26] ? 6'h1a : _ans_30_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_165 = _ans_30_leadingZeros_T_93[25] ? 6'h19 : _ans_30_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_166 = _ans_30_leadingZeros_T_93[24] ? 6'h18 : _ans_30_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_167 = _ans_30_leadingZeros_T_93[23] ? 6'h17 : _ans_30_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_168 = _ans_30_leadingZeros_T_93[22] ? 6'h16 : _ans_30_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_169 = _ans_30_leadingZeros_T_93[21] ? 6'h15 : _ans_30_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_170 = _ans_30_leadingZeros_T_93[20] ? 6'h14 : _ans_30_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_171 = _ans_30_leadingZeros_T_93[19] ? 6'h13 : _ans_30_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_172 = _ans_30_leadingZeros_T_93[18] ? 6'h12 : _ans_30_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_173 = _ans_30_leadingZeros_T_93[17] ? 6'h11 : _ans_30_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_174 = _ans_30_leadingZeros_T_93[16] ? 6'h10 : _ans_30_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_175 = _ans_30_leadingZeros_T_93[15] ? 6'hf : _ans_30_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_176 = _ans_30_leadingZeros_T_93[14] ? 6'he : _ans_30_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_177 = _ans_30_leadingZeros_T_93[13] ? 6'hd : _ans_30_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_178 = _ans_30_leadingZeros_T_93[12] ? 6'hc : _ans_30_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_179 = _ans_30_leadingZeros_T_93[11] ? 6'hb : _ans_30_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_180 = _ans_30_leadingZeros_T_93[10] ? 6'ha : _ans_30_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_181 = _ans_30_leadingZeros_T_93[9] ? 6'h9 : _ans_30_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_182 = _ans_30_leadingZeros_T_93[8] ? 6'h8 : _ans_30_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_183 = _ans_30_leadingZeros_T_93[7] ? 6'h7 : _ans_30_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_184 = _ans_30_leadingZeros_T_93[6] ? 6'h6 : _ans_30_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_185 = _ans_30_leadingZeros_T_93[5] ? 6'h5 : _ans_30_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_186 = _ans_30_leadingZeros_T_93[4] ? 6'h4 : _ans_30_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_187 = _ans_30_leadingZeros_T_93[3] ? 6'h3 : _ans_30_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_188 = _ans_30_leadingZeros_T_93[2] ? 6'h2 : _ans_30_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_leadingZeros_T_189 = _ans_30_leadingZeros_T_93[1] ? 6'h1 : _ans_30_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_30_leadingZeros = _ans_30_leadingZeros_T_93[0] ? 6'h0 : _ans_30_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_30_expRaw_T_1 = 6'h1f - ans_30_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_30_expRaw = ans_30_isZero ? 6'h0 : _ans_30_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_30_shiftAmt_T_2 = ans_30_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_30_shiftAmt = ans_30_expRaw > 6'h3 ? _ans_30_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_30_mantissaRaw_T = ans_30_absClipped >> ans_30_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_30_mantissaRaw = _ans_30_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_30_mantissa = ans_30_expRaw >= 6'h3 ? ans_30_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_30_expAdjusted = ans_30_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_30_exp_T_4 = ans_30_expAdjusted > 7'hf ? 4'hf : ans_30_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_30_exp = ans_30_isZero ? 4'h0 : _ans_30_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_30_fp8 = {ans_30_clippedX[31],ans_30_exp,ans_30_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [31:0] biasExtended_31 = {24'h0,linear_bias_31}; // @[src/main/scala/Multiple/LinearCompute.scala 150:31]
  wire [31:0] sum32_31 = tempSum_31 + biasExtended_31; // @[src/main/scala/Multiple/LinearCompute.scala 151:32]
  wire  ans_31_sign = sum32_31[31]; // @[src/main/scala/Multiple/LinearCompute.scala 31:21]
  wire [31:0] _ans_31_absX_T = ~sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 32:31]
  wire [31:0] _ans_31_absX_T_2 = _ans_31_absX_T + 32'h1; // @[src/main/scala/Multiple/LinearCompute.scala 32:34]
  wire [31:0] ans_31_absX = ans_31_sign ? _ans_31_absX_T_2 : sum32_31; // @[src/main/scala/Multiple/LinearCompute.scala 32:23]
  wire [31:0] _ans_31_shiftedX_T_1 = _GEN_14432 - ans_31_absX; // @[src/main/scala/Multiple/LinearCompute.scala 35:44]
  wire [31:0] _ans_31_shiftedX_T_3 = ans_31_absX - _GEN_14432; // @[src/main/scala/Multiple/LinearCompute.scala 35:57]
  wire [31:0] ans_31_shiftedX = ans_31_sign ? _ans_31_shiftedX_T_1 : _ans_31_shiftedX_T_3; // @[src/main/scala/Multiple/LinearCompute.scala 35:27]
  wire [48:0] _ans_31_scaledX_T_1 = ans_31_shiftedX * 17'h10000; // @[src/main/scala/Multiple/LinearCompute.scala 36:33]
  wire [48:0] ans_31_scaledX = _ans_31_scaledX_T_1 / io_scale; // @[src/main/scala/Multiple/LinearCompute.scala 36:48]
  wire [48:0] _ans_31_clippedX_T_2 = ans_31_scaledX < 49'hfffffe40 ? 49'hfffffe40 : ans_31_scaledX; // @[src/main/scala/Multiple/LinearCompute.scala 43:59]
  wire [48:0] ans_31_clippedX = ans_31_scaledX > 49'h1c0 ? 49'h1c0 : _ans_31_clippedX_T_2; // @[src/main/scala/Multiple/LinearCompute.scala 43:27]
  wire [48:0] _ans_31_absClipped_T_1 = ~ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:45]
  wire [48:0] _ans_31_absClipped_T_3 = _ans_31_absClipped_T_1 + 49'h1; // @[src/main/scala/Multiple/LinearCompute.scala 46:55]
  wire [48:0] ans_31_absClipped = ans_31_clippedX[31] ? _ans_31_absClipped_T_3 : ans_31_clippedX; // @[src/main/scala/Multiple/LinearCompute.scala 46:29]
  wire  ans_31_isZero = ans_31_absClipped == 49'h0; // @[src/main/scala/Multiple/LinearCompute.scala 47:33]
  wire [31:0] _GEN_40055 = {{16'd0}, ans_31_absClipped[31:16]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_4 = _GEN_40055 & 32'hffff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_6 = {ans_31_absClipped[15:0], 16'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_8 = _ans_31_leadingZeros_T_6 & 32'hffff0000; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_9 = _ans_31_leadingZeros_T_4 | _ans_31_leadingZeros_T_8; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40056 = {{8'd0}, _ans_31_leadingZeros_T_9[31:8]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_14 = _GEN_40056 & 32'hff00ff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_16 = {_ans_31_leadingZeros_T_9[23:0], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_18 = _ans_31_leadingZeros_T_16 & 32'hff00ff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_19 = _ans_31_leadingZeros_T_14 | _ans_31_leadingZeros_T_18; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40057 = {{4'd0}, _ans_31_leadingZeros_T_19[31:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_24 = _GEN_40057 & 32'hf0f0f0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_26 = {_ans_31_leadingZeros_T_19[27:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_28 = _ans_31_leadingZeros_T_26 & 32'hf0f0f0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_29 = _ans_31_leadingZeros_T_24 | _ans_31_leadingZeros_T_28; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40058 = {{2'd0}, _ans_31_leadingZeros_T_29[31:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_34 = _GEN_40058 & 32'h33333333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_36 = {_ans_31_leadingZeros_T_29[29:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_38 = _ans_31_leadingZeros_T_36 & 32'hcccccccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_39 = _ans_31_leadingZeros_T_34 | _ans_31_leadingZeros_T_38; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _GEN_40059 = {{1'd0}, _ans_31_leadingZeros_T_39[31:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_44 = _GEN_40059 & 32'h55555555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_46 = {_ans_31_leadingZeros_T_39[30:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_48 = _ans_31_leadingZeros_T_46 & 32'haaaaaaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [31:0] _ans_31_leadingZeros_T_49 = _ans_31_leadingZeros_T_44 | _ans_31_leadingZeros_T_48; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40060 = {{8'd0}, ans_31_absClipped[47:40]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_55 = _GEN_40060 & 16'hff; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_57 = {ans_31_absClipped[39:32], 8'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_59 = _ans_31_leadingZeros_T_57 & 16'hff00; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_60 = _ans_31_leadingZeros_T_55 | _ans_31_leadingZeros_T_59; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40061 = {{4'd0}, _ans_31_leadingZeros_T_60[15:4]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_65 = _GEN_40061 & 16'hf0f; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_67 = {_ans_31_leadingZeros_T_60[11:0], 4'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_69 = _ans_31_leadingZeros_T_67 & 16'hf0f0; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_70 = _ans_31_leadingZeros_T_65 | _ans_31_leadingZeros_T_69; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40062 = {{2'd0}, _ans_31_leadingZeros_T_70[15:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_75 = _GEN_40062 & 16'h3333; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_77 = {_ans_31_leadingZeros_T_70[13:0], 2'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_79 = _ans_31_leadingZeros_T_77 & 16'hcccc; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_80 = _ans_31_leadingZeros_T_75 | _ans_31_leadingZeros_T_79; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _GEN_40063 = {{1'd0}, _ans_31_leadingZeros_T_80[15:1]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_85 = _GEN_40063 & 16'h5555; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_87 = {_ans_31_leadingZeros_T_80[14:0], 1'h0}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_89 = _ans_31_leadingZeros_T_87 & 16'haaaa; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [15:0] _ans_31_leadingZeros_T_90 = _ans_31_leadingZeros_T_85 | _ans_31_leadingZeros_T_89; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [48:0] _ans_31_leadingZeros_T_93 = {_ans_31_leadingZeros_T_49,_ans_31_leadingZeros_T_90,ans_31_absClipped[48]}; // @[src/main/scala/Multiple/LinearCompute.scala 48:51]
  wire [5:0] _ans_31_leadingZeros_T_143 = _ans_31_leadingZeros_T_93[47] ? 6'h2f : 6'h30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_144 = _ans_31_leadingZeros_T_93[46] ? 6'h2e : _ans_31_leadingZeros_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_145 = _ans_31_leadingZeros_T_93[45] ? 6'h2d : _ans_31_leadingZeros_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_146 = _ans_31_leadingZeros_T_93[44] ? 6'h2c : _ans_31_leadingZeros_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_147 = _ans_31_leadingZeros_T_93[43] ? 6'h2b : _ans_31_leadingZeros_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_148 = _ans_31_leadingZeros_T_93[42] ? 6'h2a : _ans_31_leadingZeros_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_149 = _ans_31_leadingZeros_T_93[41] ? 6'h29 : _ans_31_leadingZeros_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_150 = _ans_31_leadingZeros_T_93[40] ? 6'h28 : _ans_31_leadingZeros_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_151 = _ans_31_leadingZeros_T_93[39] ? 6'h27 : _ans_31_leadingZeros_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_152 = _ans_31_leadingZeros_T_93[38] ? 6'h26 : _ans_31_leadingZeros_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_153 = _ans_31_leadingZeros_T_93[37] ? 6'h25 : _ans_31_leadingZeros_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_154 = _ans_31_leadingZeros_T_93[36] ? 6'h24 : _ans_31_leadingZeros_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_155 = _ans_31_leadingZeros_T_93[35] ? 6'h23 : _ans_31_leadingZeros_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_156 = _ans_31_leadingZeros_T_93[34] ? 6'h22 : _ans_31_leadingZeros_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_157 = _ans_31_leadingZeros_T_93[33] ? 6'h21 : _ans_31_leadingZeros_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_158 = _ans_31_leadingZeros_T_93[32] ? 6'h20 : _ans_31_leadingZeros_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_159 = _ans_31_leadingZeros_T_93[31] ? 6'h1f : _ans_31_leadingZeros_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_160 = _ans_31_leadingZeros_T_93[30] ? 6'h1e : _ans_31_leadingZeros_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_161 = _ans_31_leadingZeros_T_93[29] ? 6'h1d : _ans_31_leadingZeros_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_162 = _ans_31_leadingZeros_T_93[28] ? 6'h1c : _ans_31_leadingZeros_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_163 = _ans_31_leadingZeros_T_93[27] ? 6'h1b : _ans_31_leadingZeros_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_164 = _ans_31_leadingZeros_T_93[26] ? 6'h1a : _ans_31_leadingZeros_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_165 = _ans_31_leadingZeros_T_93[25] ? 6'h19 : _ans_31_leadingZeros_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_166 = _ans_31_leadingZeros_T_93[24] ? 6'h18 : _ans_31_leadingZeros_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_167 = _ans_31_leadingZeros_T_93[23] ? 6'h17 : _ans_31_leadingZeros_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_168 = _ans_31_leadingZeros_T_93[22] ? 6'h16 : _ans_31_leadingZeros_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_169 = _ans_31_leadingZeros_T_93[21] ? 6'h15 : _ans_31_leadingZeros_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_170 = _ans_31_leadingZeros_T_93[20] ? 6'h14 : _ans_31_leadingZeros_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_171 = _ans_31_leadingZeros_T_93[19] ? 6'h13 : _ans_31_leadingZeros_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_172 = _ans_31_leadingZeros_T_93[18] ? 6'h12 : _ans_31_leadingZeros_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_173 = _ans_31_leadingZeros_T_93[17] ? 6'h11 : _ans_31_leadingZeros_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_174 = _ans_31_leadingZeros_T_93[16] ? 6'h10 : _ans_31_leadingZeros_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_175 = _ans_31_leadingZeros_T_93[15] ? 6'hf : _ans_31_leadingZeros_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_176 = _ans_31_leadingZeros_T_93[14] ? 6'he : _ans_31_leadingZeros_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_177 = _ans_31_leadingZeros_T_93[13] ? 6'hd : _ans_31_leadingZeros_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_178 = _ans_31_leadingZeros_T_93[12] ? 6'hc : _ans_31_leadingZeros_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_179 = _ans_31_leadingZeros_T_93[11] ? 6'hb : _ans_31_leadingZeros_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_180 = _ans_31_leadingZeros_T_93[10] ? 6'ha : _ans_31_leadingZeros_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_181 = _ans_31_leadingZeros_T_93[9] ? 6'h9 : _ans_31_leadingZeros_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_182 = _ans_31_leadingZeros_T_93[8] ? 6'h8 : _ans_31_leadingZeros_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_183 = _ans_31_leadingZeros_T_93[7] ? 6'h7 : _ans_31_leadingZeros_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_184 = _ans_31_leadingZeros_T_93[6] ? 6'h6 : _ans_31_leadingZeros_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_185 = _ans_31_leadingZeros_T_93[5] ? 6'h5 : _ans_31_leadingZeros_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_186 = _ans_31_leadingZeros_T_93[4] ? 6'h4 : _ans_31_leadingZeros_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_187 = _ans_31_leadingZeros_T_93[3] ? 6'h3 : _ans_31_leadingZeros_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_188 = _ans_31_leadingZeros_T_93[2] ? 6'h2 : _ans_31_leadingZeros_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_leadingZeros_T_189 = _ans_31_leadingZeros_T_93[1] ? 6'h1 : _ans_31_leadingZeros_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] ans_31_leadingZeros = _ans_31_leadingZeros_T_93[0] ? 6'h0 : _ans_31_leadingZeros_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _ans_31_expRaw_T_1 = 6'h1f - ans_31_leadingZeros; // @[src/main/scala/Multiple/LinearCompute.scala 49:44]
  wire [5:0] ans_31_expRaw = ans_31_isZero ? 6'h0 : _ans_31_expRaw_T_1; // @[src/main/scala/Multiple/LinearCompute.scala 49:25]
  wire [5:0] _ans_31_shiftAmt_T_2 = ans_31_expRaw - 6'h3; // @[src/main/scala/Multiple/LinearCompute.scala 55:49]
  wire [5:0] ans_31_shiftAmt = ans_31_expRaw > 6'h3 ? _ans_31_shiftAmt_T_2 : 6'h0; // @[src/main/scala/Multiple/LinearCompute.scala 55:27]
  wire [48:0] _ans_31_mantissaRaw_T = ans_31_absClipped >> ans_31_shiftAmt; // @[src/main/scala/Multiple/LinearCompute.scala 56:39]
  wire [6:0] ans_31_mantissaRaw = _ans_31_mantissaRaw_T[6:0]; // @[src/main/scala/Multiple/LinearCompute.scala 56:51]
  wire [2:0] ans_31_mantissa = ans_31_expRaw >= 6'h3 ? ans_31_mantissaRaw[2:0] : 3'h0; // @[src/main/scala/Multiple/LinearCompute.scala 57:27]
  wire [6:0] ans_31_expAdjusted = ans_31_expRaw + 6'h7; // @[src/main/scala/Multiple/LinearCompute.scala 59:34]
  wire [3:0] _ans_31_exp_T_4 = ans_31_expAdjusted > 7'hf ? 4'hf : ans_31_expAdjusted[3:0]; // @[src/main/scala/Multiple/LinearCompute.scala 60:39]
  wire [3:0] ans_31_exp = ans_31_isZero ? 4'h0 : _ans_31_exp_T_4; // @[src/main/scala/Multiple/LinearCompute.scala 60:22]
  wire [7:0] ans_31_fp8 = {ans_31_clippedX[31],ans_31_exp,ans_31_mantissa}; // @[src/main/scala/Multiple/LinearCompute.scala 62:22]
  wire [7:0] io_featuresOut_0_scaledX = {{2'd0}, ans_0[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_0_sum = io_featuresOut_0_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_0_minVal = io_featuresOut_0_sum < 8'h40 ? io_featuresOut_0_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_1_scaledX = {{2'd0}, ans_1[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_1_sum = io_featuresOut_1_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_1_minVal = io_featuresOut_1_sum < 8'h40 ? io_featuresOut_1_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_2_scaledX = {{2'd0}, ans_2[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_2_sum = io_featuresOut_2_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_2_minVal = io_featuresOut_2_sum < 8'h40 ? io_featuresOut_2_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_3_scaledX = {{2'd0}, ans_3[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_3_sum = io_featuresOut_3_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_3_minVal = io_featuresOut_3_sum < 8'h40 ? io_featuresOut_3_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_4_scaledX = {{2'd0}, ans_4[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_4_sum = io_featuresOut_4_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_4_minVal = io_featuresOut_4_sum < 8'h40 ? io_featuresOut_4_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_5_scaledX = {{2'd0}, ans_5[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_5_sum = io_featuresOut_5_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_5_minVal = io_featuresOut_5_sum < 8'h40 ? io_featuresOut_5_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_6_scaledX = {{2'd0}, ans_6[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_6_sum = io_featuresOut_6_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_6_minVal = io_featuresOut_6_sum < 8'h40 ? io_featuresOut_6_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_7_scaledX = {{2'd0}, ans_7[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_7_sum = io_featuresOut_7_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_7_minVal = io_featuresOut_7_sum < 8'h40 ? io_featuresOut_7_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_8_scaledX = {{2'd0}, ans_8[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_8_sum = io_featuresOut_8_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_8_minVal = io_featuresOut_8_sum < 8'h40 ? io_featuresOut_8_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_9_scaledX = {{2'd0}, ans_9[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_9_sum = io_featuresOut_9_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_9_minVal = io_featuresOut_9_sum < 8'h40 ? io_featuresOut_9_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_10_scaledX = {{2'd0}, ans_10[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_10_sum = io_featuresOut_10_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_10_minVal = io_featuresOut_10_sum < 8'h40 ? io_featuresOut_10_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_11_scaledX = {{2'd0}, ans_11[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_11_sum = io_featuresOut_11_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_11_minVal = io_featuresOut_11_sum < 8'h40 ? io_featuresOut_11_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_12_scaledX = {{2'd0}, ans_12[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_12_sum = io_featuresOut_12_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_12_minVal = io_featuresOut_12_sum < 8'h40 ? io_featuresOut_12_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_13_scaledX = {{2'd0}, ans_13[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_13_sum = io_featuresOut_13_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_13_minVal = io_featuresOut_13_sum < 8'h40 ? io_featuresOut_13_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_14_scaledX = {{2'd0}, ans_14[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_14_sum = io_featuresOut_14_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_14_minVal = io_featuresOut_14_sum < 8'h40 ? io_featuresOut_14_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_15_scaledX = {{2'd0}, ans_15[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_15_sum = io_featuresOut_15_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_15_minVal = io_featuresOut_15_sum < 8'h40 ? io_featuresOut_15_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_16_scaledX = {{2'd0}, ans_16[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_16_sum = io_featuresOut_16_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_16_minVal = io_featuresOut_16_sum < 8'h40 ? io_featuresOut_16_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_17_scaledX = {{2'd0}, ans_17[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_17_sum = io_featuresOut_17_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_17_minVal = io_featuresOut_17_sum < 8'h40 ? io_featuresOut_17_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_18_scaledX = {{2'd0}, ans_18[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_18_sum = io_featuresOut_18_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_18_minVal = io_featuresOut_18_sum < 8'h40 ? io_featuresOut_18_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_19_scaledX = {{2'd0}, ans_19[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_19_sum = io_featuresOut_19_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_19_minVal = io_featuresOut_19_sum < 8'h40 ? io_featuresOut_19_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_20_scaledX = {{2'd0}, ans_20[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_20_sum = io_featuresOut_20_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_20_minVal = io_featuresOut_20_sum < 8'h40 ? io_featuresOut_20_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_21_scaledX = {{2'd0}, ans_21[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_21_sum = io_featuresOut_21_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_21_minVal = io_featuresOut_21_sum < 8'h40 ? io_featuresOut_21_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_22_scaledX = {{2'd0}, ans_22[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_22_sum = io_featuresOut_22_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_22_minVal = io_featuresOut_22_sum < 8'h40 ? io_featuresOut_22_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_23_scaledX = {{2'd0}, ans_23[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_23_sum = io_featuresOut_23_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_23_minVal = io_featuresOut_23_sum < 8'h40 ? io_featuresOut_23_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_24_scaledX = {{2'd0}, ans_24[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_24_sum = io_featuresOut_24_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_24_minVal = io_featuresOut_24_sum < 8'h40 ? io_featuresOut_24_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_25_scaledX = {{2'd0}, ans_25[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_25_sum = io_featuresOut_25_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_25_minVal = io_featuresOut_25_sum < 8'h40 ? io_featuresOut_25_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_26_scaledX = {{2'd0}, ans_26[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_26_sum = io_featuresOut_26_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_26_minVal = io_featuresOut_26_sum < 8'h40 ? io_featuresOut_26_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_27_scaledX = {{2'd0}, ans_27[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_27_sum = io_featuresOut_27_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_27_minVal = io_featuresOut_27_sum < 8'h40 ? io_featuresOut_27_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_28_scaledX = {{2'd0}, ans_28[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_28_sum = io_featuresOut_28_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_28_minVal = io_featuresOut_28_sum < 8'h40 ? io_featuresOut_28_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_29_scaledX = {{2'd0}, ans_29[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_29_sum = io_featuresOut_29_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_29_minVal = io_featuresOut_29_sum < 8'h40 ? io_featuresOut_29_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_30_scaledX = {{2'd0}, ans_30[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_30_sum = io_featuresOut_30_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_30_minVal = io_featuresOut_30_sum < 8'h40 ? io_featuresOut_30_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  wire [7:0] io_featuresOut_31_scaledX = {{2'd0}, ans_31[7:2]}; // @[src/main/scala/Multiple/LinearCompute.scala 159:27 160:17]
  wire [7:0] io_featuresOut_31_sum = io_featuresOut_31_scaledX + 8'h20; // @[src/main/scala/Multiple/LinearCompute.scala 162:24]
  wire [7:0] io_featuresOut_31_minVal = io_featuresOut_31_sum < 8'h40 ? io_featuresOut_31_sum : 8'h40; // @[src/main/scala/Multiple/LinearCompute.scala 164:25]
  reg  regs__0; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__1; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__2; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg  regs__3; // @[src/main/scala/fpga/Pipeline.scala 41:31]
  reg [2047:0] regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  reg [2047:0] regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 32:31]
  assign io_pipe_validOut = regs__3; // @[src/main/scala/fpga/Pipeline.scala 46:21]
  assign io_pipe_phvOut = regs_1_3; // @[src/main/scala/fpga/Pipeline.scala 37:21]
  assign io_featuresOut_0 = io_featuresOut_0_minVal > 8'h0 ? io_featuresOut_0_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_1 = io_featuresOut_1_minVal > 8'h0 ? io_featuresOut_1_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_2 = io_featuresOut_2_minVal > 8'h0 ? io_featuresOut_2_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_3 = io_featuresOut_3_minVal > 8'h0 ? io_featuresOut_3_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_4 = io_featuresOut_4_minVal > 8'h0 ? io_featuresOut_4_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_5 = io_featuresOut_5_minVal > 8'h0 ? io_featuresOut_5_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_6 = io_featuresOut_6_minVal > 8'h0 ? io_featuresOut_6_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_7 = io_featuresOut_7_minVal > 8'h0 ? io_featuresOut_7_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_8 = io_featuresOut_8_minVal > 8'h0 ? io_featuresOut_8_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_9 = io_featuresOut_9_minVal > 8'h0 ? io_featuresOut_9_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_10 = io_featuresOut_10_minVal > 8'h0 ? io_featuresOut_10_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_11 = io_featuresOut_11_minVal > 8'h0 ? io_featuresOut_11_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_12 = io_featuresOut_12_minVal > 8'h0 ? io_featuresOut_12_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_13 = io_featuresOut_13_minVal > 8'h0 ? io_featuresOut_13_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_14 = io_featuresOut_14_minVal > 8'h0 ? io_featuresOut_14_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_15 = io_featuresOut_15_minVal > 8'h0 ? io_featuresOut_15_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_16 = io_featuresOut_16_minVal > 8'h0 ? io_featuresOut_16_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_17 = io_featuresOut_17_minVal > 8'h0 ? io_featuresOut_17_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_18 = io_featuresOut_18_minVal > 8'h0 ? io_featuresOut_18_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_19 = io_featuresOut_19_minVal > 8'h0 ? io_featuresOut_19_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_20 = io_featuresOut_20_minVal > 8'h0 ? io_featuresOut_20_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_21 = io_featuresOut_21_minVal > 8'h0 ? io_featuresOut_21_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_22 = io_featuresOut_22_minVal > 8'h0 ? io_featuresOut_22_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_23 = io_featuresOut_23_minVal > 8'h0 ? io_featuresOut_23_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_24 = io_featuresOut_24_minVal > 8'h0 ? io_featuresOut_24_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_25 = io_featuresOut_25_minVal > 8'h0 ? io_featuresOut_25_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_26 = io_featuresOut_26_minVal > 8'h0 ? io_featuresOut_26_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_27 = io_featuresOut_27_minVal > 8'h0 ? io_featuresOut_27_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_28 = io_featuresOut_28_minVal > 8'h0 ? io_featuresOut_28_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_29 = io_featuresOut_29_minVal > 8'h0 ? io_featuresOut_29_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_30 = io_featuresOut_30_minVal > 8'h0 ? io_featuresOut_30_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  assign io_featuresOut_31 = io_featuresOut_31_minVal > 8'h0 ? io_featuresOut_31_minVal : 8'h0; // @[src/main/scala/Multiple/LinearCompute.scala 165:25]
  always @(posedge clock) begin
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h0 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_0 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_1 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h2 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_2 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h3 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_3 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h4 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_4 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h5 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_5 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h6 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_6 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h7 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_7 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h8 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_8 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h9 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_9 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'ha == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_10 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'hb == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_11 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'hc == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_12 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'hd == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_13 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'he == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_14 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'hf == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_15 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h10 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_16 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h11 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_17 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h12 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_18 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h13 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_19 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h14 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_20 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h15 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_21 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h16 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_22 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h17 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_23 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h18 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_24 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h19 == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_25 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1a == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_26 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1b == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_27 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1c == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_28 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1d == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_29 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1e == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_30 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (io_config_weight) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (6'h3f == io_config_i[5:0] & 5'h1f == io_config_j[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
          linear_weight_63_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 23:53]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h0 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_0 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_1 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h2 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_2 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h3 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_3 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h4 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_4 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h5 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_5 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h6 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_6 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h7 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_7 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h8 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_8 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h9 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_9 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'ha == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_10 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'hb == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_11 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'hc == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_12 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'hd == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_13 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'he == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_14 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'hf == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_15 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h10 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_16 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h11 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_17 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h12 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_18 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h13 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_19 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h14 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_20 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h15 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_21 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h16 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_22 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h17 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_23 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h18 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_24 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h19 == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_25 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1a == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_26 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1b == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_27 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1c == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_28 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1d == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_29 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1e == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_30 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (io_config_en) begin // @[src/main/scala/Multiple/LinearCompute.scala 21:25]
      if (!(io_config_weight)) begin // @[src/main/scala/Multiple/LinearCompute.scala 22:33]
        if (5'h1f == io_config_i[4:0]) begin // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
          linear_bias_31 <= io_config_value; // @[src/main/scala/Multiple/LinearCompute.scala 25:38]
        end
      end
    end
    if (weightQ8_63_0_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_0 <= 8'h0;
    end else begin
      weightQ8_63_0 <= weightQ8_63_0_fp8;
    end
    if (weightQ8_63_1_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_1 <= 8'h0;
    end else begin
      weightQ8_63_1 <= weightQ8_63_1_fp8;
    end
    if (weightQ8_63_2_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_2 <= 8'h0;
    end else begin
      weightQ8_63_2 <= weightQ8_63_2_fp8;
    end
    if (weightQ8_63_3_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_3 <= 8'h0;
    end else begin
      weightQ8_63_3 <= weightQ8_63_3_fp8;
    end
    if (weightQ8_63_4_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_4 <= 8'h0;
    end else begin
      weightQ8_63_4 <= weightQ8_63_4_fp8;
    end
    if (weightQ8_63_5_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_5 <= 8'h0;
    end else begin
      weightQ8_63_5 <= weightQ8_63_5_fp8;
    end
    if (weightQ8_63_6_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_6 <= 8'h0;
    end else begin
      weightQ8_63_6 <= weightQ8_63_6_fp8;
    end
    if (weightQ8_63_7_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_7 <= 8'h0;
    end else begin
      weightQ8_63_7 <= weightQ8_63_7_fp8;
    end
    if (weightQ8_63_8_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_8 <= 8'h0;
    end else begin
      weightQ8_63_8 <= weightQ8_63_8_fp8;
    end
    if (weightQ8_63_9_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_9 <= 8'h0;
    end else begin
      weightQ8_63_9 <= weightQ8_63_9_fp8;
    end
    if (weightQ8_63_10_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_10 <= 8'h0;
    end else begin
      weightQ8_63_10 <= weightQ8_63_10_fp8;
    end
    if (weightQ8_63_11_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_11 <= 8'h0;
    end else begin
      weightQ8_63_11 <= weightQ8_63_11_fp8;
    end
    if (weightQ8_63_12_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_12 <= 8'h0;
    end else begin
      weightQ8_63_12 <= weightQ8_63_12_fp8;
    end
    if (weightQ8_63_13_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_13 <= 8'h0;
    end else begin
      weightQ8_63_13 <= weightQ8_63_13_fp8;
    end
    if (weightQ8_63_14_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_14 <= 8'h0;
    end else begin
      weightQ8_63_14 <= weightQ8_63_14_fp8;
    end
    if (weightQ8_63_15_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_15 <= 8'h0;
    end else begin
      weightQ8_63_15 <= weightQ8_63_15_fp8;
    end
    if (weightQ8_63_16_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_16 <= 8'h0;
    end else begin
      weightQ8_63_16 <= weightQ8_63_16_fp8;
    end
    if (weightQ8_63_17_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_17 <= 8'h0;
    end else begin
      weightQ8_63_17 <= weightQ8_63_17_fp8;
    end
    if (weightQ8_63_18_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_18 <= 8'h0;
    end else begin
      weightQ8_63_18 <= weightQ8_63_18_fp8;
    end
    if (weightQ8_63_19_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_19 <= 8'h0;
    end else begin
      weightQ8_63_19 <= weightQ8_63_19_fp8;
    end
    if (weightQ8_63_20_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_20 <= 8'h0;
    end else begin
      weightQ8_63_20 <= weightQ8_63_20_fp8;
    end
    if (weightQ8_63_21_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_21 <= 8'h0;
    end else begin
      weightQ8_63_21 <= weightQ8_63_21_fp8;
    end
    if (weightQ8_63_22_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_22 <= 8'h0;
    end else begin
      weightQ8_63_22 <= weightQ8_63_22_fp8;
    end
    if (weightQ8_63_23_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_23 <= 8'h0;
    end else begin
      weightQ8_63_23 <= weightQ8_63_23_fp8;
    end
    if (weightQ8_63_24_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_24 <= 8'h0;
    end else begin
      weightQ8_63_24 <= weightQ8_63_24_fp8;
    end
    if (weightQ8_63_25_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_25 <= 8'h0;
    end else begin
      weightQ8_63_25 <= weightQ8_63_25_fp8;
    end
    if (weightQ8_63_26_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_26 <= 8'h0;
    end else begin
      weightQ8_63_26 <= weightQ8_63_26_fp8;
    end
    if (weightQ8_63_27_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_27 <= 8'h0;
    end else begin
      weightQ8_63_27 <= weightQ8_63_27_fp8;
    end
    if (weightQ8_63_28_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_28 <= 8'h0;
    end else begin
      weightQ8_63_28 <= weightQ8_63_28_fp8;
    end
    if (weightQ8_63_29_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_29 <= 8'h0;
    end else begin
      weightQ8_63_29 <= weightQ8_63_29_fp8;
    end
    if (weightQ8_63_30_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_30 <= 8'h0;
    end else begin
      weightQ8_63_30 <= weightQ8_63_30_fp8;
    end
    if (weightQ8_63_31_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      weightQ8_63_31 <= 8'h0;
    end else begin
      weightQ8_63_31 <= weightQ8_63_31_fp8;
    end
    if (ansAll_63_0_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_0 <= _ansAll_63_0_T_4;
    end else begin
      ansAll_63_0 <= ansAll_63_0_resultAbs;
    end
    if (ansAll_63_1_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_1 <= _ansAll_63_1_T_4;
    end else begin
      ansAll_63_1 <= ansAll_63_1_resultAbs;
    end
    if (ansAll_63_2_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_2 <= _ansAll_63_2_T_4;
    end else begin
      ansAll_63_2 <= ansAll_63_2_resultAbs;
    end
    if (ansAll_63_3_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_3 <= _ansAll_63_3_T_4;
    end else begin
      ansAll_63_3 <= ansAll_63_3_resultAbs;
    end
    if (ansAll_63_4_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_4 <= _ansAll_63_4_T_4;
    end else begin
      ansAll_63_4 <= ansAll_63_4_resultAbs;
    end
    if (ansAll_63_5_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_5 <= _ansAll_63_5_T_4;
    end else begin
      ansAll_63_5 <= ansAll_63_5_resultAbs;
    end
    if (ansAll_63_6_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_6 <= _ansAll_63_6_T_4;
    end else begin
      ansAll_63_6 <= ansAll_63_6_resultAbs;
    end
    if (ansAll_63_7_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_7 <= _ansAll_63_7_T_4;
    end else begin
      ansAll_63_7 <= ansAll_63_7_resultAbs;
    end
    if (ansAll_63_8_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_8 <= _ansAll_63_8_T_4;
    end else begin
      ansAll_63_8 <= ansAll_63_8_resultAbs;
    end
    if (ansAll_63_9_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_9 <= _ansAll_63_9_T_4;
    end else begin
      ansAll_63_9 <= ansAll_63_9_resultAbs;
    end
    if (ansAll_63_10_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_10 <= _ansAll_63_10_T_4;
    end else begin
      ansAll_63_10 <= ansAll_63_10_resultAbs;
    end
    if (ansAll_63_11_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_11 <= _ansAll_63_11_T_4;
    end else begin
      ansAll_63_11 <= ansAll_63_11_resultAbs;
    end
    if (ansAll_63_12_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_12 <= _ansAll_63_12_T_4;
    end else begin
      ansAll_63_12 <= ansAll_63_12_resultAbs;
    end
    if (ansAll_63_13_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_13 <= _ansAll_63_13_T_4;
    end else begin
      ansAll_63_13 <= ansAll_63_13_resultAbs;
    end
    if (ansAll_63_14_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_14 <= _ansAll_63_14_T_4;
    end else begin
      ansAll_63_14 <= ansAll_63_14_resultAbs;
    end
    if (ansAll_63_15_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_15 <= _ansAll_63_15_T_4;
    end else begin
      ansAll_63_15 <= ansAll_63_15_resultAbs;
    end
    if (ansAll_63_16_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_16 <= _ansAll_63_16_T_4;
    end else begin
      ansAll_63_16 <= ansAll_63_16_resultAbs;
    end
    if (ansAll_63_17_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_17 <= _ansAll_63_17_T_4;
    end else begin
      ansAll_63_17 <= ansAll_63_17_resultAbs;
    end
    if (ansAll_63_18_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_18 <= _ansAll_63_18_T_4;
    end else begin
      ansAll_63_18 <= ansAll_63_18_resultAbs;
    end
    if (ansAll_63_19_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_19 <= _ansAll_63_19_T_4;
    end else begin
      ansAll_63_19 <= ansAll_63_19_resultAbs;
    end
    if (ansAll_63_20_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_20 <= _ansAll_63_20_T_4;
    end else begin
      ansAll_63_20 <= ansAll_63_20_resultAbs;
    end
    if (ansAll_63_21_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_21 <= _ansAll_63_21_T_4;
    end else begin
      ansAll_63_21 <= ansAll_63_21_resultAbs;
    end
    if (ansAll_63_22_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_22 <= _ansAll_63_22_T_4;
    end else begin
      ansAll_63_22 <= ansAll_63_22_resultAbs;
    end
    if (ansAll_63_23_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_23 <= _ansAll_63_23_T_4;
    end else begin
      ansAll_63_23 <= ansAll_63_23_resultAbs;
    end
    if (ansAll_63_24_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_24 <= _ansAll_63_24_T_4;
    end else begin
      ansAll_63_24 <= ansAll_63_24_resultAbs;
    end
    if (ansAll_63_25_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_25 <= _ansAll_63_25_T_4;
    end else begin
      ansAll_63_25 <= ansAll_63_25_resultAbs;
    end
    if (ansAll_63_26_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_26 <= _ansAll_63_26_T_4;
    end else begin
      ansAll_63_26 <= ansAll_63_26_resultAbs;
    end
    if (ansAll_63_27_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_27 <= _ansAll_63_27_T_4;
    end else begin
      ansAll_63_27 <= ansAll_63_27_resultAbs;
    end
    if (ansAll_63_28_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_28 <= _ansAll_63_28_T_4;
    end else begin
      ansAll_63_28 <= ansAll_63_28_resultAbs;
    end
    if (ansAll_63_29_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_29 <= _ansAll_63_29_T_4;
    end else begin
      ansAll_63_29 <= ansAll_63_29_resultAbs;
    end
    if (ansAll_63_30_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_30 <= _ansAll_63_30_T_4;
    end else begin
      ansAll_63_30 <= ansAll_63_30_resultAbs;
    end
    if (ansAll_63_31_signProd) begin // @[src/main/scala/Multiple/LinearCompute.scala 110:12]
      ansAll_63_31 <= _ansAll_63_31_T_4;
    end else begin
      ansAll_63_31 <= ansAll_63_31_resultAbs;
    end
    if (ans_0_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_0 <= 8'h0;
    end else begin
      ans_0 <= ans_0_fp8;
    end
    if (ans_1_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_1 <= 8'h0;
    end else begin
      ans_1 <= ans_1_fp8;
    end
    if (ans_2_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_2 <= 8'h0;
    end else begin
      ans_2 <= ans_2_fp8;
    end
    if (ans_3_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_3 <= 8'h0;
    end else begin
      ans_3 <= ans_3_fp8;
    end
    if (ans_4_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_4 <= 8'h0;
    end else begin
      ans_4 <= ans_4_fp8;
    end
    if (ans_5_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_5 <= 8'h0;
    end else begin
      ans_5 <= ans_5_fp8;
    end
    if (ans_6_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_6 <= 8'h0;
    end else begin
      ans_6 <= ans_6_fp8;
    end
    if (ans_7_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_7 <= 8'h0;
    end else begin
      ans_7 <= ans_7_fp8;
    end
    if (ans_8_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_8 <= 8'h0;
    end else begin
      ans_8 <= ans_8_fp8;
    end
    if (ans_9_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_9 <= 8'h0;
    end else begin
      ans_9 <= ans_9_fp8;
    end
    if (ans_10_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_10 <= 8'h0;
    end else begin
      ans_10 <= ans_10_fp8;
    end
    if (ans_11_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_11 <= 8'h0;
    end else begin
      ans_11 <= ans_11_fp8;
    end
    if (ans_12_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_12 <= 8'h0;
    end else begin
      ans_12 <= ans_12_fp8;
    end
    if (ans_13_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_13 <= 8'h0;
    end else begin
      ans_13 <= ans_13_fp8;
    end
    if (ans_14_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_14 <= 8'h0;
    end else begin
      ans_14 <= ans_14_fp8;
    end
    if (ans_15_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_15 <= 8'h0;
    end else begin
      ans_15 <= ans_15_fp8;
    end
    if (ans_16_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_16 <= 8'h0;
    end else begin
      ans_16 <= ans_16_fp8;
    end
    if (ans_17_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_17 <= 8'h0;
    end else begin
      ans_17 <= ans_17_fp8;
    end
    if (ans_18_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_18 <= 8'h0;
    end else begin
      ans_18 <= ans_18_fp8;
    end
    if (ans_19_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_19 <= 8'h0;
    end else begin
      ans_19 <= ans_19_fp8;
    end
    if (ans_20_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_20 <= 8'h0;
    end else begin
      ans_20 <= ans_20_fp8;
    end
    if (ans_21_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_21 <= 8'h0;
    end else begin
      ans_21 <= ans_21_fp8;
    end
    if (ans_22_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_22 <= 8'h0;
    end else begin
      ans_22 <= ans_22_fp8;
    end
    if (ans_23_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_23 <= 8'h0;
    end else begin
      ans_23 <= ans_23_fp8;
    end
    if (ans_24_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_24 <= 8'h0;
    end else begin
      ans_24 <= ans_24_fp8;
    end
    if (ans_25_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_25 <= 8'h0;
    end else begin
      ans_25 <= ans_25_fp8;
    end
    if (ans_26_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_26 <= 8'h0;
    end else begin
      ans_26 <= ans_26_fp8;
    end
    if (ans_27_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_27 <= 8'h0;
    end else begin
      ans_27 <= ans_27_fp8;
    end
    if (ans_28_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_28 <= 8'h0;
    end else begin
      ans_28 <= ans_28_fp8;
    end
    if (ans_29_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_29 <= 8'h0;
    end else begin
      ans_29 <= ans_29_fp8;
    end
    if (ans_30_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_30 <= 8'h0;
    end else begin
      ans_30 <= ans_30_fp8;
    end
    if (ans_31_isZero) begin // @[src/main/scala/Multiple/LinearCompute.scala 63:12]
      ans_31 <= 8'h0;
    end else begin
      ans_31 <= ans_31_fp8;
    end
    tempSum_0 <= tempSum_0 + ansAll_63_0; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_1 <= tempSum_1 + ansAll_63_1; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_2 <= tempSum_2 + ansAll_63_2; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_3 <= tempSum_3 + ansAll_63_3; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_4 <= tempSum_4 + ansAll_63_4; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_5 <= tempSum_5 + ansAll_63_5; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_6 <= tempSum_6 + ansAll_63_6; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_7 <= tempSum_7 + ansAll_63_7; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_8 <= tempSum_8 + ansAll_63_8; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_9 <= tempSum_9 + ansAll_63_9; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_10 <= tempSum_10 + ansAll_63_10; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_11 <= tempSum_11 + ansAll_63_11; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_12 <= tempSum_12 + ansAll_63_12; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_13 <= tempSum_13 + ansAll_63_13; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_14 <= tempSum_14 + ansAll_63_14; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_15 <= tempSum_15 + ansAll_63_15; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_16 <= tempSum_16 + ansAll_63_16; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_17 <= tempSum_17 + ansAll_63_17; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_18 <= tempSum_18 + ansAll_63_18; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_19 <= tempSum_19 + ansAll_63_19; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_20 <= tempSum_20 + ansAll_63_20; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_21 <= tempSum_21 + ansAll_63_21; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_22 <= tempSum_22 + ansAll_63_22; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_23 <= tempSum_23 + ansAll_63_23; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_24 <= tempSum_24 + ansAll_63_24; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_25 <= tempSum_25 + ansAll_63_25; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_26 <= tempSum_26 + ansAll_63_26; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_27 <= tempSum_27 + ansAll_63_27; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_28 <= tempSum_28 + ansAll_63_28; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_29 <= tempSum_29 + ansAll_63_29; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_30 <= tempSum_30 + ansAll_63_30; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    tempSum_31 <= tempSum_31 + ansAll_63_31; // @[src/main/scala/Multiple/LinearCompute.scala 144:38]
    regs__0 <= io_pipe_validIn; // @[src/main/scala/fpga/Pipeline.scala 45:25]
    regs__1 <= regs__0; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__2 <= regs__1; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs__3 <= regs__2; // @[src/main/scala/fpga/Pipeline.scala 43:37]
    regs_1_0 <= io_pipe_phvIn; // @[src/main/scala/fpga/Pipeline.scala 36:25]
    regs_1_1 <= regs_1_0; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_2 <= regs_1_1; // @[src/main/scala/fpga/Pipeline.scala 34:37]
    regs_1_3 <= regs_1_2; // @[src/main/scala/fpga/Pipeline.scala 34:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  linear_weight_63_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  linear_weight_63_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  linear_weight_63_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  linear_weight_63_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  linear_weight_63_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  linear_weight_63_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  linear_weight_63_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  linear_weight_63_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  linear_weight_63_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  linear_weight_63_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  linear_weight_63_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  linear_weight_63_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  linear_weight_63_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  linear_weight_63_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  linear_weight_63_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  linear_weight_63_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  linear_weight_63_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  linear_weight_63_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  linear_weight_63_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  linear_weight_63_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  linear_weight_63_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  linear_weight_63_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  linear_weight_63_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  linear_weight_63_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  linear_weight_63_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  linear_weight_63_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  linear_weight_63_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  linear_weight_63_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  linear_weight_63_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  linear_weight_63_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  linear_weight_63_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  linear_weight_63_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  linear_bias_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  linear_bias_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  linear_bias_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  linear_bias_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  linear_bias_4 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  linear_bias_5 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  linear_bias_6 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  linear_bias_7 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  linear_bias_8 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  linear_bias_9 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  linear_bias_10 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  linear_bias_11 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  linear_bias_12 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  linear_bias_13 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  linear_bias_14 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  linear_bias_15 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  linear_bias_16 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  linear_bias_17 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  linear_bias_18 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  linear_bias_19 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  linear_bias_20 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  linear_bias_21 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  linear_bias_22 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  linear_bias_23 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  linear_bias_24 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  linear_bias_25 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  linear_bias_26 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  linear_bias_27 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  linear_bias_28 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  linear_bias_29 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  linear_bias_30 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  linear_bias_31 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  weightQ8_63_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  weightQ8_63_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  weightQ8_63_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  weightQ8_63_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  weightQ8_63_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  weightQ8_63_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  weightQ8_63_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  weightQ8_63_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  weightQ8_63_8 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  weightQ8_63_9 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  weightQ8_63_10 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  weightQ8_63_11 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  weightQ8_63_12 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  weightQ8_63_13 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  weightQ8_63_14 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  weightQ8_63_15 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  weightQ8_63_16 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  weightQ8_63_17 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  weightQ8_63_18 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  weightQ8_63_19 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  weightQ8_63_20 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  weightQ8_63_21 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  weightQ8_63_22 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  weightQ8_63_23 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  weightQ8_63_24 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  weightQ8_63_25 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  weightQ8_63_26 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  weightQ8_63_27 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  weightQ8_63_28 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  weightQ8_63_29 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  weightQ8_63_30 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  weightQ8_63_31 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  ansAll_63_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  ansAll_63_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  ansAll_63_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  ansAll_63_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  ansAll_63_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  ansAll_63_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  ansAll_63_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  ansAll_63_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  ansAll_63_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  ansAll_63_9 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  ansAll_63_10 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  ansAll_63_11 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  ansAll_63_12 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  ansAll_63_13 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  ansAll_63_14 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  ansAll_63_15 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  ansAll_63_16 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  ansAll_63_17 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  ansAll_63_18 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  ansAll_63_19 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  ansAll_63_20 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  ansAll_63_21 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  ansAll_63_22 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  ansAll_63_23 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  ansAll_63_24 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  ansAll_63_25 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  ansAll_63_26 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  ansAll_63_27 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  ansAll_63_28 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  ansAll_63_29 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  ansAll_63_30 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  ansAll_63_31 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  ans_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  ans_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  ans_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  ans_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  ans_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  ans_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  ans_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  ans_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  ans_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  ans_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  ans_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  ans_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  ans_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  ans_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  ans_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  ans_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  ans_16 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  ans_17 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  ans_18 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  ans_19 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  ans_20 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  ans_21 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  ans_22 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  ans_23 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  ans_24 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  ans_25 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  ans_26 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  ans_27 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  ans_28 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  ans_29 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  ans_30 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  ans_31 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  tempSum_0 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  tempSum_1 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  tempSum_2 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  tempSum_3 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  tempSum_4 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  tempSum_5 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  tempSum_6 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  tempSum_7 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  tempSum_8 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  tempSum_9 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  tempSum_10 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  tempSum_11 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  tempSum_12 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  tempSum_13 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  tempSum_14 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  tempSum_15 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  tempSum_16 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  tempSum_17 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  tempSum_18 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  tempSum_19 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  tempSum_20 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  tempSum_21 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  tempSum_22 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  tempSum_23 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  tempSum_24 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  tempSum_25 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  tempSum_26 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  tempSum_27 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  tempSum_28 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  tempSum_29 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  tempSum_30 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  tempSum_31 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  regs__0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  regs__1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  regs__2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  regs__3 = _RAND_195[0:0];
  _RAND_196 = {64{`RANDOM}};
  regs_1_0 = _RAND_196[2047:0];
  _RAND_197 = {64{`RANDOM}};
  regs_1_1 = _RAND_197[2047:0];
  _RAND_198 = {64{`RANDOM}};
  regs_1_2 = _RAND_198[2047:0];
  _RAND_199 = {64{`RANDOM}};
  regs_1_3 = _RAND_199[2047:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
