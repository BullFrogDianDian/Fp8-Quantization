module FloatMul8(
  input        clock,
  input        reset,
  input  [7:0] io_a, // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 7:16]
  input  [7:0] io_b, // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 7:16]
  output [7:0] io_c // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 7:16]
);
  wire  a_sign = io_a[7]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 20:22]
  wire [3:0] a_exp = io_a[6:3]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 21:21]
  wire [2:0] a_mant = io_a[2:0]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 22:22]
  wire  b_sign = io_b[7]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 24:22]
  wire [3:0] b_exp = io_b[6:3]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 25:21]
  wire [2:0] b_mant = io_b[2:0]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 26:22]
  wire  res_sign = a_sign ^ b_sign; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 29:27]
  wire [3:0] a_mant_full = {1'h1,a_mant}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 32:26]
  wire [3:0] b_mant_full = {1'h1,b_mant}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 33:26]
  wire [7:0] mant_product = a_mant_full * b_mant_full; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 36:36]
  wire  normalize = mant_product[7]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 39:33]
  wire [2:0] norm_mant = normalize ? mant_product[6:4] : mant_product[5:3]; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 40:24]
  wire [4:0] exp_sum = a_exp + b_exp; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 43:25]
  wire [5:0] _res_exp_T = exp_sum - 5'h7; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 44:27]
  wire [5:0] _GEN_4 = {{5'd0}, normalize}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 44:34]
  wire [5:0] res_exp = _res_exp_T + _GEN_4; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 44:34]
  wire  a_zero = a_exp == 4'h0; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 47:24]
  wire  b_zero = b_exp == 4'h0; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 48:24]
  wire  a_inf = a_exp == 4'hf; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 49:23]
  wire  b_inf = b_exp == 4'hf; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 50:23]
  wire [7:0] _result_T = {res_sign,7'h0}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 57:22]
  wire [7:0] _result_T_1 = {res_sign,4'hf,3'h0}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 60:22]
  wire [7:0] _result_T_5 = {res_sign,res_exp[3:0],norm_mant}; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 69:22]
  wire [7:0] _GEN_0 = res_exp == 6'h0 | res_exp[4] ? _result_T : _result_T_5; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 64:47 66:16 69:16]
  wire [7:0] _GEN_1 = res_exp >= 6'hf ? _result_T_1 : _GEN_0; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 61:33 63:16]
  wire [7:0] _GEN_2 = a_inf | b_inf ? _result_T_1 : _GEN_1; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 58:32 60:16]
  assign io_c = a_zero | b_zero ? _result_T : _GEN_2; // @[Users/apple/Desktop/floatedpoint8-1/src/main/scala/Multiple/FloatMul8.scala 55:28 57:16]
endmodule
